library ieee;
                use ieee.std_logic_1164.all;
                use ieee.numeric_std.all;
                use ieee.std_logic_unsigned.all;
                entity multiple_tests is
                end multiple_tests;
                architecture projecttb of multiple_tests is
                constant c_CLOCK_PERIOD		: time := 100 ns;
                signal   tb_done		: std_logic;
                signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
                signal   tb_rst	                : std_logic := '0';
                signal   tb_start		: std_logic := '0';
                signal   tb_clk		        : std_logic := '0';
                signal   mem_o_data,mem_i_data	: std_logic_vector (7 downto 0);
                signal   enable_wire  		: std_logic;
                signal   mem_we		        : std_logic;
                type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
                signal RAM: ram_type := (0 => "11110011",
1 => std_logic_vector(to_unsigned( 210, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 72, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 212, 8)),
10 => std_logic_vector(to_unsigned( 77, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 95, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
signal count : integer := 0;
-- MASK_OUT: 	 11110011
 component project_reti_logiche is
                port (
                    i_clk         : in  std_logic;
                    i_start       : in  std_logic;
                    i_rst         : in  std_logic;
                    i_data        : in  std_logic_vector(7 downto 0);
                    o_address     : out std_logic_vector(15 downto 0);
                    o_done        : out std_logic;
                    o_en          : out std_logic;
                    o_we          : out std_logic;
                    o_data        : out std_logic_vector (7 downto 0)
                    );
                end component project_reti_logiche;
                begin
                UUT: project_reti_logiche
                port map (
                        i_clk      	=> tb_clk,
                        i_start       => tb_start,
                        i_rst      	=> tb_rst,
                        i_data    	=> mem_o_data,
                        o_address  	=> mem_address,
                        o_done      	=> tb_done,
                        o_en   	=> enable_wire,
                        o_we 		=> mem_we,
                        o_data    	=> mem_i_data
                        );
                p_CLK_GEN : process is
                begin
                    wait for c_CLOCK_PERIOD/2;
                    tb_clk <= not tb_clk;
                end process p_CLK_GEN;
                MEM : process(tb_clk)
                begin
                    if tb_clk'event and tb_clk = '1' then
                        if enable_wire = '1' then
                            if mem_we = '1' then
                                RAM(conv_integer(mem_address))  <= mem_i_data;
                                mem_o_data                      <= mem_i_data after 2 ns;
                            else
                                mem_o_data <= RAM(conv_integer(mem_address)) after 2 ns;
                            end if;
                        end if;
                    elsif tb_rst = '1' then 
 if (count=0) then count <= 1;elsif count = 1 then count <= 2; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 90, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 25, 8)),
6 => std_logic_vector(to_unsigned( 127, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 214, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 2 then count <= 3; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 98, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 209, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 3 then count <= 4; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 96, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 217, 8)),
5 => std_logic_vector(to_unsigned( 7, 8)),
6 => std_logic_vector(to_unsigned( 200, 8)),
7 => std_logic_vector(to_unsigned( 203, 8)),
8 => std_logic_vector(to_unsigned( 10, 8)),
9 => std_logic_vector(to_unsigned( 238, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 74, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 4 then count <= 5; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 215, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 198, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 159, 8)),
9 => std_logic_vector(to_unsigned( 86, 8)),
10 => std_logic_vector(to_unsigned( 112, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 47, 8)),
14 => std_logic_vector(to_unsigned( 177, 8)),
15 => std_logic_vector(to_unsigned( 68, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 5 then count <= 6; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 171, 8)),
2 => std_logic_vector(to_unsigned( 62, 8)),
3 => std_logic_vector(to_unsigned( 218, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 203, 8)),
8 => std_logic_vector(to_unsigned( 15, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 165, 8)),
11 => std_logic_vector(to_unsigned( 255, 8)),
12 => std_logic_vector(to_unsigned( 219, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 168, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 6 then count <= 7; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 168, 8)),
13 => std_logic_vector(to_unsigned( 236, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 7 then count <= 8; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 46, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 46, 8)),
8 => std_logic_vector(to_unsigned( 127, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 75, 8)),
11 => std_logic_vector(to_unsigned( 248, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 77, 8)),
17 => std_logic_vector(to_unsigned( 46, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 8 then count <= 9; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 3, 8)),
6 => std_logic_vector(to_unsigned( 245, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 188, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 238, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 243, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 252, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 193, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 9 then count <= 10; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 245, 8)),
7 => std_logic_vector(to_unsigned( 229, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 110, 8)),
10 => std_logic_vector(to_unsigned( 210, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 245, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 201, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 10 then count <= 11; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 222, 8)),
3 => std_logic_vector(to_unsigned( 56, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 60, 8)),
8 => std_logic_vector(to_unsigned( 241, 8)),
9 => std_logic_vector(to_unsigned( 58, 8)),
10 => std_logic_vector(to_unsigned( 83, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 233, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 0, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 243, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 204, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 11 then count <= 12; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 49, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 83, 8)),
4 => std_logic_vector(to_unsigned( 75, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 21, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 138, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 213, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 12 then count <= 13; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 43, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 26, 8)),
4 => std_logic_vector(to_unsigned( 165, 8)),
5 => std_logic_vector(to_unsigned( 25, 8)),
6 => std_logic_vector(to_unsigned( 190, 8)),
7 => std_logic_vector(to_unsigned( 13, 8)),
8 => std_logic_vector(to_unsigned( 249, 8)),
9 => std_logic_vector(to_unsigned( 23, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 78, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 29, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 44, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 13 then count <= 14; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 102, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 251, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 209, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 64, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 14 then count <= 15; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 237, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 249, 8)),
6 => std_logic_vector(to_unsigned( 32, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 15, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 77, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 126, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 15 then count <= 16; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 28, 8)),
2 => std_logic_vector(to_unsigned( 142, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 190, 8)),
6 => std_logic_vector(to_unsigned( 193, 8)),
7 => std_logic_vector(to_unsigned( 223, 8)),
8 => std_logic_vector(to_unsigned( 131, 8)),
9 => std_logic_vector(to_unsigned( 57, 8)),
10 => std_logic_vector(to_unsigned( 180, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 191, 8)),
13 => std_logic_vector(to_unsigned( 44, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110010
elsif count = 16 then count <= 17; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 19, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 149, 8)),
9 => std_logic_vector(to_unsigned( 148, 8)),
10 => std_logic_vector(to_unsigned( 155, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 17 then count <= 18; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 196, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 209, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 207, 8)),
8 => std_logic_vector(to_unsigned( 205, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 217, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 31, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 199, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00010111
elsif count = 18 then count <= 19; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 54, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 181, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 168, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011001
elsif count = 19 then count <= 20; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 140, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 166, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 107, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 66, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 242, 8)),
16 => std_logic_vector(to_unsigned( 54, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 20 then count <= 21; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 239, 8)),
2 => std_logic_vector(to_unsigned( 13, 8)),
3 => std_logic_vector(to_unsigned( 41, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 236, 8)),
7 => std_logic_vector(to_unsigned( 98, 8)),
8 => std_logic_vector(to_unsigned( 34, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 27, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 138, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 44, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 21 then count <= 22; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 42, 8)),
2 => std_logic_vector(to_unsigned( 153, 8)),
3 => std_logic_vector(to_unsigned( 237, 8)),
4 => std_logic_vector(to_unsigned( 237, 8)),
5 => std_logic_vector(to_unsigned( 249, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 200, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 41, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 87, 8)),
14 => std_logic_vector(to_unsigned( 80, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 22 then count <= 23; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 130, 8)),
2 => std_logic_vector(to_unsigned( 201, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 245, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 221, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 229, 8)),
14 => std_logic_vector(to_unsigned( 172, 8)),
15 => std_logic_vector(to_unsigned( 63, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 23 then count <= 24; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 83, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 197, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 202, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 221, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 226, 8)),
15 => std_logic_vector(to_unsigned( 51, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 56, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 24 then count <= 25; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 37, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 241, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 75, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 17, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 25 then count <= 26; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 242, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 179, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 74, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 203, 8)),
15 => std_logic_vector(to_unsigned( 227, 8)),
16 => std_logic_vector(to_unsigned( 29, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 26 then count <= 27; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 253, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 240, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 117, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 206, 8)),
13 => std_logic_vector(to_unsigned( 6, 8)),
14 => std_logic_vector(to_unsigned( 234, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 27 then count <= 28; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 45, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 122, 8)),
6 => std_logic_vector(to_unsigned( 34, 8)),
7 => std_logic_vector(to_unsigned( 161, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 146, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 17, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 28 then count <= 29; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 2, 8)),
3 => std_logic_vector(to_unsigned( 235, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 82, 8)),
6 => std_logic_vector(to_unsigned( 173, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 30, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 8, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 54, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 29 then count <= 30; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 165, 8)),
2 => std_logic_vector(to_unsigned( 118, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 90, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 154, 8)),
14 => std_logic_vector(to_unsigned( 146, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 30 then count <= 31; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 141, 8)),
3 => std_logic_vector(to_unsigned( 4, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 12, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 141, 8)),
8 => std_logic_vector(to_unsigned( 182, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 238, 8)),
11 => std_logic_vector(to_unsigned( 163, 8)),
12 => std_logic_vector(to_unsigned( 18, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 206, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 31 then count <= 32; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 214, 8)),
4 => std_logic_vector(to_unsigned( 77, 8)),
5 => std_logic_vector(to_unsigned( 217, 8)),
6 => std_logic_vector(to_unsigned( 80, 8)),
7 => std_logic_vector(to_unsigned( 188, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 250, 8)),
11 => std_logic_vector(to_unsigned( 207, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 213, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 32 then count <= 33; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 46, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 177, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 28, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 103, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 33 then count <= 34; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 129, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 180, 8)),
8 => std_logic_vector(to_unsigned( 22, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 237, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 25, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 49, 8)),
17 => std_logic_vector(to_unsigned( 184, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 34 then count <= 35; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 94, 8)),
3 => std_logic_vector(to_unsigned( 181, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 161, 8)),
6 => std_logic_vector(to_unsigned( 19, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 59, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 3, 8)),
12 => std_logic_vector(to_unsigned( 57, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 167, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 35 then count <= 36; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 13, 8)),
4 => std_logic_vector(to_unsigned( 199, 8)),
5 => std_logic_vector(to_unsigned( 215, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 217, 8)),
8 => std_logic_vector(to_unsigned( 46, 8)),
9 => std_logic_vector(to_unsigned( 176, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 218, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 211, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 172, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 36 then count <= 37; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 120, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 116, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 16, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 213, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00001111
elsif count = 37 then count <= 38; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 44, 8)),
2 => std_logic_vector(to_unsigned( 28, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 205, 8)),
6 => std_logic_vector(to_unsigned( 59, 8)),
7 => std_logic_vector(to_unsigned( 223, 8)),
8 => std_logic_vector(to_unsigned( 77, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 2, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 52, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 38 then count <= 39; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 216, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 108, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 108, 8)),
8 => std_logic_vector(to_unsigned( 57, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 129, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 41, 8)),
15 => std_logic_vector(to_unsigned( 103, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 39 then count <= 40; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 195, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 146, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 24, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 40, 8)),
16 => std_logic_vector(to_unsigned( 214, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 40 then count <= 41; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 213, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 66, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 83, 8)),
11 => std_logic_vector(to_unsigned( 1, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 3, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 204, 8)),
18 => std_logic_vector(to_unsigned( 63, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011001
elsif count = 41 then count <= 42; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 91, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 47, 8)),
5 => std_logic_vector(to_unsigned( 85, 8)),
6 => std_logic_vector(to_unsigned( 44, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 100, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 12, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 42 then count <= 43; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 233, 8)),
3 => std_logic_vector(to_unsigned( 75, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 225, 8)),
13 => std_logic_vector(to_unsigned( 7, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 17, 8)),
16 => std_logic_vector(to_unsigned( 231, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 197, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 43 then count <= 44; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 48, 8)),
4 => std_logic_vector(to_unsigned( 54, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 28, 8)),
8 => std_logic_vector(to_unsigned( 32, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 56, 8)),
11 => std_logic_vector(to_unsigned( 233, 8)),
12 => std_logic_vector(to_unsigned( 145, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 47, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 251, 8)),
17 => std_logic_vector(to_unsigned( 61, 8)),
18 => std_logic_vector(to_unsigned( 33, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 44 then count <= 45; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 223, 8)),
2 => std_logic_vector(to_unsigned( 40, 8)),
3 => std_logic_vector(to_unsigned( 181, 8)),
4 => std_logic_vector(to_unsigned( 72, 8)),
5 => std_logic_vector(to_unsigned( 213, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 236, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 213, 8)),
13 => std_logic_vector(to_unsigned( 214, 8)),
14 => std_logic_vector(to_unsigned( 31, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 14, 8)),
17 => std_logic_vector(to_unsigned( 204, 8)),
18 => std_logic_vector(to_unsigned( 58, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 45 then count <= 46; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 182, 8)),
3 => std_logic_vector(to_unsigned( 14, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 73, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 13, 8)),
11 => std_logic_vector(to_unsigned( 191, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 45, 8)),
15 => std_logic_vector(to_unsigned( 209, 8)),
16 => std_logic_vector(to_unsigned( 183, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 48, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 46 then count <= 47; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 232, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 161, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 116, 8)),
8 => std_logic_vector(to_unsigned( 97, 8)),
9 => std_logic_vector(to_unsigned( 81, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 38, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 251, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 47 then count <= 48; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 64, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 56, 8)),
9 => std_logic_vector(to_unsigned( 63, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 244, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 47, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 48 then count <= 49; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 235, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 171, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 23, 8)),
6 => std_logic_vector(to_unsigned( 249, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 236, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 241, 8)),
14 => std_logic_vector(to_unsigned( 52, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 249, 8)),
17 => std_logic_vector(to_unsigned( 197, 8)),
18 => std_logic_vector(to_unsigned( 48, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 49 then count <= 50; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 27, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 31, 8)),
9 => std_logic_vector(to_unsigned( 222, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 51, 8)),
13 => std_logic_vector(to_unsigned( 154, 8)),
14 => std_logic_vector(to_unsigned( 90, 8)),
15 => std_logic_vector(to_unsigned( 143, 8)),
16 => std_logic_vector(to_unsigned( 79, 8)),
17 => std_logic_vector(to_unsigned( 196, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 50 then count <= 51; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 91, 8)),
2 => std_logic_vector(to_unsigned( 212, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 203, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 240, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 211, 8)),
9 => std_logic_vector(to_unsigned( 107, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 51, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 209, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010011
elsif count = 51 then count <= 52; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 81, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 226, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 83, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 52 then count <= 53; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 123, 8)),
5 => std_logic_vector(to_unsigned( 142, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 183, 8)),
8 => std_logic_vector(to_unsigned( 191, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 137, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 39, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 213, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010111
elsif count = 53 then count <= 54; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 212, 8)),
2 => std_logic_vector(to_unsigned( 26, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 1, 8)),
6 => std_logic_vector(to_unsigned( 192, 8)),
7 => std_logic_vector(to_unsigned( 213, 8)),
8 => std_logic_vector(to_unsigned( 27, 8)),
9 => std_logic_vector(to_unsigned( 177, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 54, 8)),
13 => std_logic_vector(to_unsigned( 233, 8)),
14 => std_logic_vector(to_unsigned( 253, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 197, 8)),
18 => std_logic_vector(to_unsigned( 46, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 54 then count <= 55; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 136, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 63, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 54, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 78, 8)),
13 => std_logic_vector(to_unsigned( 229, 8)),
14 => std_logic_vector(to_unsigned( 228, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 8, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00100111
elsif count = 55 then count <= 56; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 59, 8)),
2 => std_logic_vector(to_unsigned( 247, 8)),
3 => std_logic_vector(to_unsigned( 254, 8)),
4 => std_logic_vector(to_unsigned( 226, 8)),
5 => std_logic_vector(to_unsigned( 98, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 119, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 203, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 56 then count <= 57; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 95, 8)),
5 => std_logic_vector(to_unsigned( 82, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 46, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 191, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 73, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 174, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 57 then count <= 58; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 40, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 111, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 191, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 58 then count <= 59; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 92, 8)),
2 => std_logic_vector(to_unsigned( 125, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 28, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 31, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 15, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 73, 8)),
14 => std_logic_vector(to_unsigned( 163, 8)),
15 => std_logic_vector(to_unsigned( 216, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 47, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 59 then count <= 60; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 68, 8)),
2 => std_logic_vector(to_unsigned( 201, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 207, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 37, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 22, 8)),
10 => std_logic_vector(to_unsigned( 163, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 64, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 60 then count <= 61; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 95, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 174, 8)),
8 => std_logic_vector(to_unsigned( 100, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 250, 8)),
14 => std_logic_vector(to_unsigned( 1, 8)),
15 => std_logic_vector(to_unsigned( 3, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 61 then count <= 62; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 230, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 63, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 169, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 241, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 62 then count <= 63; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 92, 8)),
2 => std_logic_vector(to_unsigned( 200, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 164, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 101, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 9, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 63 then count <= 64; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 116, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 234, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 220, 8)),
9 => std_logic_vector(to_unsigned( 130, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 191, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 108, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 64 then count <= 65; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 242, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 178, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 64, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 206, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 252, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 212, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 65 then count <= 66; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 70, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 204, 8)),
15 => std_logic_vector(to_unsigned( 198, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 66 then count <= 67; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 99, 8)),
2 => std_logic_vector(to_unsigned( 248, 8)),
3 => std_logic_vector(to_unsigned( 149, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 41, 8)),
6 => std_logic_vector(to_unsigned( 13, 8)),
7 => std_logic_vector(to_unsigned( 101, 8)),
8 => std_logic_vector(to_unsigned( 250, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 241, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 67 then count <= 68; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 4, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 30, 8)),
6 => std_logic_vector(to_unsigned( 227, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 40, 8)),
14 => std_logic_vector(to_unsigned( 254, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 54, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011010
elsif count = 68 then count <= 69; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 43, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 172, 8)),
7 => std_logic_vector(to_unsigned( 189, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 183, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 69 then count <= 70; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 230, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 53, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 238, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 70 then count <= 71; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 38, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 31, 8)),
7 => std_logic_vector(to_unsigned( 168, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 197, 8)),
14 => std_logic_vector(to_unsigned( 47, 8)),
15 => std_logic_vector(to_unsigned( 206, 8)),
16 => std_logic_vector(to_unsigned( 78, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 71 then count <= 72; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 199, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 193, 8)),
6 => std_logic_vector(to_unsigned( 142, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 218, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 211, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 190, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 241, 8)),
16 => std_logic_vector(to_unsigned( 11, 8)),
17 => std_logic_vector(to_unsigned( 200, 8)),
18 => std_logic_vector(to_unsigned( 181, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 72 then count <= 73; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 72, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 106, 8)),
5 => std_logic_vector(to_unsigned( 53, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 137, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 156, 8)),
11 => std_logic_vector(to_unsigned( 54, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 26, 8)),
14 => std_logic_vector(to_unsigned( 180, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 73 then count <= 74; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 160, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 53, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 83, 8)),
7 => std_logic_vector(to_unsigned( 238, 8)),
8 => std_logic_vector(to_unsigned( 144, 8)),
9 => std_logic_vector(to_unsigned( 217, 8)),
10 => std_logic_vector(to_unsigned( 89, 8)),
11 => std_logic_vector(to_unsigned( 190, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 90, 8)),
16 => std_logic_vector(to_unsigned( 29, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 74 then count <= 75; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 156, 8)),
6 => std_logic_vector(to_unsigned( 87, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 1, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 75 then count <= 76; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 59, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 210, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 32, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 45, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010011
elsif count = 76 then count <= 77; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 101, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 104, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 198, 8)),
8 => std_logic_vector(to_unsigned( 37, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 111, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 77 then count <= 78; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 38, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 175, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 53, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 78 then count <= 79; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 246, 8)),
4 => std_logic_vector(to_unsigned( 245, 8)),
5 => std_logic_vector(to_unsigned( 241, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 184, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 228, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 34, 8)),
13 => std_logic_vector(to_unsigned( 183, 8)),
14 => std_logic_vector(to_unsigned( 218, 8)),
15 => std_logic_vector(to_unsigned( 167, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 200, 8)),
18 => std_logic_vector(to_unsigned( 51, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 79 then count <= 80; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 130, 8)),
3 => std_logic_vector(to_unsigned( 162, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 227, 8)),
8 => std_logic_vector(to_unsigned( 23, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 49, 8)),
12 => std_logic_vector(to_unsigned( 187, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 236, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 80 then count <= 81; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 92, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 114, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 91, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 212, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 81 then count <= 82; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 32, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 141, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 79, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 233, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 224, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 82 then count <= 83; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 63, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 204, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 197, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 83 then count <= 84; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 238, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 56, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 124, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 110, 8)),
13 => std_logic_vector(to_unsigned( 71, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 84 then count <= 85; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 106, 8)),
5 => std_logic_vector(to_unsigned( 22, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 21, 8)),
8 => std_logic_vector(to_unsigned( 201, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 136, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 104, 8)),
16 => std_logic_vector(to_unsigned( 64, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 85 then count <= 86; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 202, 8)),
2 => std_logic_vector(to_unsigned( 226, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 215, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 221, 8)),
9 => std_logic_vector(to_unsigned( 156, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 215, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 67, 8)),
15 => std_logic_vector(to_unsigned( 131, 8)),
16 => std_logic_vector(to_unsigned( 63, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 86 then count <= 87; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 189, 8)),
7 => std_logic_vector(to_unsigned( 23, 8)),
8 => std_logic_vector(to_unsigned( 245, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 117, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 87 then count <= 88; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 190, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 207, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 200, 8)),
16 => std_logic_vector(to_unsigned( 56, 8)),
17 => std_logic_vector(to_unsigned( 188, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 88 then count <= 89; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 247, 8)),
2 => std_logic_vector(to_unsigned( 222, 8)),
3 => std_logic_vector(to_unsigned( 162, 8)),
4 => std_logic_vector(to_unsigned( 10, 8)),
5 => std_logic_vector(to_unsigned( 100, 8)),
6 => std_logic_vector(to_unsigned( 10, 8)),
7 => std_logic_vector(to_unsigned( 2, 8)),
8 => std_logic_vector(to_unsigned( 170, 8)),
9 => std_logic_vector(to_unsigned( 126, 8)),
10 => std_logic_vector(to_unsigned( 14, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 3, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 59, 8)),
15 => std_logic_vector(to_unsigned( 42, 8)),
16 => std_logic_vector(to_unsigned( 68, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 89 then count <= 90; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 250, 8)),
10 => std_logic_vector(to_unsigned( 0, 8)),
11 => std_logic_vector(to_unsigned( 173, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 138, 8)),
15 => std_logic_vector(to_unsigned( 4, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 90 then count <= 91; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 225, 8)),
2 => std_logic_vector(to_unsigned( 7, 8)),
3 => std_logic_vector(to_unsigned( 98, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 128, 8)),
8 => std_logic_vector(to_unsigned( 61, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 44, 8)),
11 => std_logic_vector(to_unsigned( 40, 8)),
12 => std_logic_vector(to_unsigned( 245, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 130, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 91 then count <= 92; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 36, 8)),
4 => std_logic_vector(to_unsigned( 252, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 57, 8)),
8 => std_logic_vector(to_unsigned( 245, 8)),
9 => std_logic_vector(to_unsigned( 31, 8)),
10 => std_logic_vector(to_unsigned( 239, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 131, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 163, 8)),
15 => std_logic_vector(to_unsigned( 50, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 47, 8)),
18 => std_logic_vector(to_unsigned( 208, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 92 then count <= 93; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 205, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 78, 8)),
5 => std_logic_vector(to_unsigned( 208, 8)),
6 => std_logic_vector(to_unsigned( 79, 8)),
7 => std_logic_vector(to_unsigned( 71, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 60, 8)),
12 => std_logic_vector(to_unsigned( 42, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 21, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 33, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 93 then count <= 94; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 92, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 41, 8)),
4 => std_logic_vector(to_unsigned( 71, 8)),
5 => std_logic_vector(to_unsigned( 223, 8)),
6 => std_logic_vector(to_unsigned( 185, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 198, 8)),
10 => std_logic_vector(to_unsigned( 250, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 88, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 79, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 94 then count <= 95; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 204, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 254, 8)),
13 => std_logic_vector(to_unsigned( 235, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 164, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 95 then count <= 96; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 31, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 189, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 159, 8)),
9 => std_logic_vector(to_unsigned( 25, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 211, 8)),
14 => std_logic_vector(to_unsigned( 44, 8)),
15 => std_logic_vector(to_unsigned( 152, 8)),
16 => std_logic_vector(to_unsigned( 141, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 96 then count <= 97; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 154, 8)),
4 => std_logic_vector(to_unsigned( 80, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 89, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001110
elsif count = 97 then count <= 98; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 2, 8)),
3 => std_logic_vector(to_unsigned( 28, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 31, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 224, 8)),
13 => std_logic_vector(to_unsigned( 222, 8)),
14 => std_logic_vector(to_unsigned( 13, 8)),
15 => std_logic_vector(to_unsigned( 213, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 98 then count <= 99; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 239, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 148, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 69, 8)),
9 => std_logic_vector(to_unsigned( 248, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 235, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 20, 8)),
17 => std_logic_vector(to_unsigned( 189, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 99 then count <= 100; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 49, 8)),
2 => std_logic_vector(to_unsigned( 82, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 166, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 213, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001100
elsif count = 100 then count <= 101; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 241, 8)),
2 => std_logic_vector(to_unsigned( 29, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 140, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 13, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 101 then count <= 102; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 206, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 124, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 103, 8)),
8 => std_logic_vector(to_unsigned( 144, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 25, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 102 then count <= 103; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 0, 8)),
2 => std_logic_vector(to_unsigned( 190, 8)),
3 => std_logic_vector(to_unsigned( 89, 8)),
4 => std_logic_vector(to_unsigned( 23, 8)),
5 => std_logic_vector(to_unsigned( 134, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 106, 8)),
9 => std_logic_vector(to_unsigned( 255, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 43, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 6, 8)),
14 => std_logic_vector(to_unsigned( 254, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 103 then count <= 104; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 19, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 21, 8)),
4 => std_logic_vector(to_unsigned( 55, 8)),
5 => std_logic_vector(to_unsigned( 161, 8)),
6 => std_logic_vector(to_unsigned( 7, 8)),
7 => std_logic_vector(to_unsigned( 14, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 51, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 252, 8)),
15 => std_logic_vector(to_unsigned( 7, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 81, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 104 then count <= 105; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 233, 8)),
4 => std_logic_vector(to_unsigned( 90, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 156, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 41, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 242, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 58, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 198, 8)),
16 => std_logic_vector(to_unsigned( 9, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 105 then count <= 106; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 198, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 202, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 186, 8)),
10 => std_logic_vector(to_unsigned( 177, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 99, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 106 then count <= 107; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 195, 8)),
2 => std_logic_vector(to_unsigned( 158, 8)),
3 => std_logic_vector(to_unsigned( 221, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 250, 8)),
12 => std_logic_vector(to_unsigned( 62, 8)),
13 => std_logic_vector(to_unsigned( 196, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 212, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 182, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001101
elsif count = 107 then count <= 108; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 152, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 0, 8)),
6 => std_logic_vector(to_unsigned( 160, 8)),
7 => std_logic_vector(to_unsigned( 242, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 144, 8)),
15 => std_logic_vector(to_unsigned( 194, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 108 then count <= 109; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 34, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 33, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 71, 8)),
8 => std_logic_vector(to_unsigned( 202, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 244, 8)),
14 => std_logic_vector(to_unsigned( 10, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 106, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 109 then count <= 110; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 72, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 230, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 13, 8)),
8 => std_logic_vector(to_unsigned( 22, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 163, 8)),
12 => std_logic_vector(to_unsigned( 131, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 174, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 110 then count <= 111; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 189, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 71, 8)),
11 => std_logic_vector(to_unsigned( 210, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 3, 8)),
16 => std_logic_vector(to_unsigned( 250, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 111 then count <= 112; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 193, 8)),
4 => std_logic_vector(to_unsigned( 16, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 225, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 50, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 58, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 112 then count <= 113; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 139, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 34, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 248, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 141, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 113 then count <= 114; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 237, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 214, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 22, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 233, 8)),
12 => std_logic_vector(to_unsigned( 145, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 159, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 114 then count <= 115; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 197, 8)),
2 => std_logic_vector(to_unsigned( 229, 8)),
3 => std_logic_vector(to_unsigned( 68, 8)),
4 => std_logic_vector(to_unsigned( 17, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 166, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 76, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 7, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 225, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 115 then count <= 116; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 137, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 218, 8)),
10 => std_logic_vector(to_unsigned( 183, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 24, 8)),
13 => std_logic_vector(to_unsigned( 59, 8)),
14 => std_logic_vector(to_unsigned( 214, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 116 then count <= 117; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 129, 8)),
2 => std_logic_vector(to_unsigned( 72, 8)),
3 => std_logic_vector(to_unsigned( 205, 8)),
4 => std_logic_vector(to_unsigned( 72, 8)),
5 => std_logic_vector(to_unsigned( 27, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 117, 8)),
11 => std_logic_vector(to_unsigned( 62, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 83, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 117 then count <= 118; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 227, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 33, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 165, 8)),
11 => std_logic_vector(to_unsigned( 120, 8)),
12 => std_logic_vector(to_unsigned( 228, 8)),
13 => std_logic_vector(to_unsigned( 87, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110000
elsif count = 118 then count <= 119; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 17, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 195, 8)),
5 => std_logic_vector(to_unsigned( 14, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 57, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 58, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 219, 8)),
13 => std_logic_vector(to_unsigned( 71, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 225, 8)),
17 => std_logic_vector(to_unsigned( 39, 8)),
18 => std_logic_vector(to_unsigned( 212, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 119 then count <= 120; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 41, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 98, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 216, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 188, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 158, 8)),
15 => std_logic_vector(to_unsigned( 155, 8)),
16 => std_logic_vector(to_unsigned( 214, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 183, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 120 then count <= 121; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 230, 8)),
3 => std_logic_vector(to_unsigned( 247, 8)),
4 => std_logic_vector(to_unsigned( 217, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 91, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 20, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 255, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001101
elsif count = 121 then count <= 122; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 49, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 36, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 250, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 32, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 173, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 190, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 122 then count <= 123; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 228, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 231, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 218, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 73, 8)),
14 => std_logic_vector(to_unsigned( 218, 8)),
15 => std_logic_vector(to_unsigned( 81, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00001111
elsif count = 123 then count <= 124; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 219, 8)),
4 => std_logic_vector(to_unsigned( 28, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 5, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 131, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 63, 8)),
11 => std_logic_vector(to_unsigned( 190, 8)),
12 => std_logic_vector(to_unsigned( 79, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 185, 8)),
15 => std_logic_vector(to_unsigned( 239, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 124 then count <= 125; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 45, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 67, 8)),
4 => std_logic_vector(to_unsigned( 56, 8)),
5 => std_logic_vector(to_unsigned( 77, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 33, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 74, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 60, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 125 then count <= 126; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 53, 8)),
3 => std_logic_vector(to_unsigned( 38, 8)),
4 => std_logic_vector(to_unsigned( 116, 8)),
5 => std_logic_vector(to_unsigned( 24, 8)),
6 => std_logic_vector(to_unsigned( 249, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 31, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 60, 8)),
12 => std_logic_vector(to_unsigned( 138, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 126 then count <= 127; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 98, 8)),
4 => std_logic_vector(to_unsigned( 221, 8)),
5 => std_logic_vector(to_unsigned( 20, 8)),
6 => std_logic_vector(to_unsigned( 4, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 225, 8)),
14 => std_logic_vector(to_unsigned( 73, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 193, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 181, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 127 then count <= 128; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 252, 8)),
2 => std_logic_vector(to_unsigned( 88, 8)),
3 => std_logic_vector(to_unsigned( 109, 8)),
4 => std_logic_vector(to_unsigned( 26, 8)),
5 => std_logic_vector(to_unsigned( 207, 8)),
6 => std_logic_vector(to_unsigned( 39, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 206, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 35, 8)),
11 => std_logic_vector(to_unsigned( 100, 8)),
12 => std_logic_vector(to_unsigned( 35, 8)),
13 => std_logic_vector(to_unsigned( 64, 8)),
14 => std_logic_vector(to_unsigned( 181, 8)),
15 => std_logic_vector(to_unsigned( 182, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110010
elsif count = 128 then count <= 129; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 0, 8)),
12 => std_logic_vector(to_unsigned( 179, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 129 then count <= 130; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 151, 8)),
3 => std_logic_vector(to_unsigned( 109, 8)),
4 => std_logic_vector(to_unsigned( 4, 8)),
5 => std_logic_vector(to_unsigned( 250, 8)),
6 => std_logic_vector(to_unsigned( 223, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 238, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 33, 8)),
15 => std_logic_vector(to_unsigned( 232, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 203, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 130 then count <= 131; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 5, 8)),
2 => std_logic_vector(to_unsigned( 76, 8)),
3 => std_logic_vector(to_unsigned( 17, 8)),
4 => std_logic_vector(to_unsigned( 224, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 119, 8)),
13 => std_logic_vector(to_unsigned( 163, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 162, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 131 then count <= 132; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 26, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 164, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 247, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 8, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 132 then count <= 133; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 74, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 21, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 56, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 133 then count <= 134; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 8, 8)),
2 => std_logic_vector(to_unsigned( 241, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 193, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 44, 8)),
13 => std_logic_vector(to_unsigned( 253, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 52, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 134 then count <= 135; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 161, 8)),
6 => std_logic_vector(to_unsigned( 45, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 197, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 238, 8)),
16 => std_logic_vector(to_unsigned( 10, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 135 then count <= 136; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 34, 8)),
2 => std_logic_vector(to_unsigned( 60, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 215, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 174, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 80, 8)),
10 => std_logic_vector(to_unsigned( 205, 8)),
11 => std_logic_vector(to_unsigned( 111, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 140, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 103, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 136 then count <= 137; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 83, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 47, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 172, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 114, 8)),
10 => std_logic_vector(to_unsigned( 255, 8)),
11 => std_logic_vector(to_unsigned( 38, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 74, 8)),
14 => std_logic_vector(to_unsigned( 69, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 137 then count <= 138; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 225, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 196, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 242, 8)),
14 => std_logic_vector(to_unsigned( 244, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 138 then count <= 139; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 199, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 227, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 251, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 196, 8)),
14 => std_logic_vector(to_unsigned( 146, 8)),
15 => std_logic_vector(to_unsigned( 185, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 186, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001101
elsif count = 139 then count <= 140; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 28, 8)),
3 => std_logic_vector(to_unsigned( 159, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 132, 8)),
10 => std_logic_vector(to_unsigned( 234, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 1, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 181, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 133, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001110
elsif count = 140 then count <= 141; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 149, 8)),
6 => std_logic_vector(to_unsigned( 95, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 31, 8)),
9 => std_logic_vector(to_unsigned( 232, 8)),
10 => std_logic_vector(to_unsigned( 4, 8)),
11 => std_logic_vector(to_unsigned( 131, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 24, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 51, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 141 then count <= 142; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 239, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 142 then count <= 143; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 39, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 32, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 215, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 223, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 43, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 31, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00001111
elsif count = 143 then count <= 144; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 140, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 68, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 204, 8)),
10 => std_logic_vector(to_unsigned( 44, 8)),
11 => std_logic_vector(to_unsigned( 226, 8)),
12 => std_logic_vector(to_unsigned( 244, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 75, 8)),
15 => std_logic_vector(to_unsigned( 92, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 144 then count <= 145; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 92, 8)),
2 => std_logic_vector(to_unsigned( 209, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 42, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 225, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 173, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 239, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 5, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 202, 8)),
17 => std_logic_vector(to_unsigned( 73, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 145 then count <= 146; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 79, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 70, 8)),
4 => std_logic_vector(to_unsigned( 41, 8)),
5 => std_logic_vector(to_unsigned( 58, 8)),
6 => std_logic_vector(to_unsigned( 53, 8)),
7 => std_logic_vector(to_unsigned( 209, 8)),
8 => std_logic_vector(to_unsigned( 6, 8)),
9 => std_logic_vector(to_unsigned( 110, 8)),
10 => std_logic_vector(to_unsigned( 89, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 247, 8)),
13 => std_logic_vector(to_unsigned( 105, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 51, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010111
elsif count = 146 then count <= 147; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 182, 8)),
4 => std_logic_vector(to_unsigned( 41, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 240, 8)),
7 => std_logic_vector(to_unsigned( 10, 8)),
8 => std_logic_vector(to_unsigned( 179, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 37, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 80, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 147 then count <= 148; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 240, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 227, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 1, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 188, 8)),
12 => std_logic_vector(to_unsigned( 84, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 170, 8)),
17 => std_logic_vector(to_unsigned( 188, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 148 then count <= 149; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 165, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 166, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 201, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 23, 8)),
13 => std_logic_vector(to_unsigned( 217, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 92, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 128, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 149 then count <= 150; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 171, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 24, 8)),
6 => std_logic_vector(to_unsigned( 148, 8)),
7 => std_logic_vector(to_unsigned( 94, 8)),
8 => std_logic_vector(to_unsigned( 23, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 89, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 150 then count <= 151; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 178, 8)),
4 => std_logic_vector(to_unsigned( 227, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 229, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 155, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 147, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 80, 8)),
15 => std_logic_vector(to_unsigned( 185, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 151 then count <= 152; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 215, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 170, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 116, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 0, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 152 then count <= 153; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 60, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 221, 8)),
5 => std_logic_vector(to_unsigned( 131, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 227, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 182, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 153 then count <= 154; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 79, 8)),
4 => std_logic_vector(to_unsigned( 232, 8)),
5 => std_logic_vector(to_unsigned( 124, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 23, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 68, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 154 then count <= 155; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 209, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 238, 8)),
14 => std_logic_vector(to_unsigned( 158, 8)),
15 => std_logic_vector(to_unsigned( 252, 8)),
16 => std_logic_vector(to_unsigned( 54, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 155 then count <= 156; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 248, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 119, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 86, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 131, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 156 then count <= 157; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 171, 8)),
2 => std_logic_vector(to_unsigned( 230, 8)),
3 => std_logic_vector(to_unsigned( 224, 8)),
4 => std_logic_vector(to_unsigned( 66, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 133, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 113, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 157 then count <= 158; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 182, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 97, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 107, 8)),
12 => std_logic_vector(to_unsigned( 50, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 252, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 158 then count <= 159; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 78, 8)),
2 => std_logic_vector(to_unsigned( 28, 8)),
3 => std_logic_vector(to_unsigned( 81, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 218, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 45, 8)),
12 => std_logic_vector(to_unsigned( 61, 8)),
13 => std_logic_vector(to_unsigned( 252, 8)),
14 => std_logic_vector(to_unsigned( 246, 8)),
15 => std_logic_vector(to_unsigned( 173, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 159 then count <= 160; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 211, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 212, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 216, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 242, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00010111
elsif count = 160 then count <= 161; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 233, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 213, 8)),
7 => std_logic_vector(to_unsigned( 240, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 181, 8)),
15 => std_logic_vector(to_unsigned( 204, 8)),
16 => std_logic_vector(to_unsigned( 26, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 161 then count <= 162; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 195, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 207, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 172, 8)),
13 => std_logic_vector(to_unsigned( 209, 8)),
14 => std_logic_vector(to_unsigned( 179, 8)),
15 => std_logic_vector(to_unsigned( 233, 8)),
16 => std_logic_vector(to_unsigned( 105, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 162 then count <= 163; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 36, 8)),
4 => std_logic_vector(to_unsigned( 204, 8)),
5 => std_logic_vector(to_unsigned( 208, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 188, 8)),
10 => std_logic_vector(to_unsigned( 29, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 247, 8)),
13 => std_logic_vector(to_unsigned( 249, 8)),
14 => std_logic_vector(to_unsigned( 255, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001101
elsif count = 163 then count <= 164; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 230, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 89, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 53, 8)),
14 => std_logic_vector(to_unsigned( 37, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 207, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 164 then count <= 165; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 16, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 161, 8)),
6 => std_logic_vector(to_unsigned( 53, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 4, 8)),
9 => std_logic_vector(to_unsigned( 182, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 26, 8)),
13 => std_logic_vector(to_unsigned( 173, 8)),
14 => std_logic_vector(to_unsigned( 35, 8)),
15 => std_logic_vector(to_unsigned( 177, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 206, 8)),
18 => std_logic_vector(to_unsigned( 50, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 165 then count <= 166; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 153, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 101, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 29, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 206, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 166 then count <= 167; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 95, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 4, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 202, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 87, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 71, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 35, 8)),
16 => std_logic_vector(to_unsigned( 98, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 167 then count <= 168; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 30, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 67, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 243, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 251, 8)),
11 => std_logic_vector(to_unsigned( 240, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 51, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 37, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 168 then count <= 169; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 227, 8)),
2 => std_logic_vector(to_unsigned( 3, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 197, 8)),
11 => std_logic_vector(to_unsigned( 206, 8)),
12 => std_logic_vector(to_unsigned( 235, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 181, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 169 then count <= 170; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 93, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 184, 8)),
8 => std_logic_vector(to_unsigned( 46, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 8, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 46, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 170 then count <= 171; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 163, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 216, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 169, 8)),
9 => std_logic_vector(to_unsigned( 216, 8)),
10 => std_logic_vector(to_unsigned( 10, 8)),
11 => std_logic_vector(to_unsigned( 204, 8)),
12 => std_logic_vector(to_unsigned( 179, 8)),
13 => std_logic_vector(to_unsigned( 225, 8)),
14 => std_logic_vector(to_unsigned( 158, 8)),
15 => std_logic_vector(to_unsigned( 170, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 149, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 171 then count <= 172; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 212, 8)),
6 => std_logic_vector(to_unsigned( 3, 8)),
7 => std_logic_vector(to_unsigned( 199, 8)),
8 => std_logic_vector(to_unsigned( 55, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 203, 8)),
12 => std_logic_vector(to_unsigned( 59, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 25, 8)),
17 => std_logic_vector(to_unsigned( 219, 8)),
18 => std_logic_vector(to_unsigned( 44, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 172 then count <= 173; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 141, 8)),
2 => std_logic_vector(to_unsigned( 36, 8)),
3 => std_logic_vector(to_unsigned( 250, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 24, 8)),
6 => std_logic_vector(to_unsigned( 89, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 104, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 118, 8)),
18 => std_logic_vector(to_unsigned( 54, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 173 then count <= 174; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 255, 8)),
2 => std_logic_vector(to_unsigned( 32, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 251, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 183, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 254, 8)),
12 => std_logic_vector(to_unsigned( 10, 8)),
13 => std_logic_vector(to_unsigned( 236, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 211, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 174 then count <= 175; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 110, 8)),
10 => std_logic_vector(to_unsigned( 237, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 244, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 175 then count <= 176; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 50, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 15, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 52, 8)),
13 => std_logic_vector(to_unsigned( 71, 8)),
14 => std_logic_vector(to_unsigned( 141, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 176 then count <= 177; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 204, 8)),
5 => std_logic_vector(to_unsigned( 204, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 249, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 253, 8)),
13 => std_logic_vector(to_unsigned( 218, 8)),
14 => std_logic_vector(to_unsigned( 144, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 182, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010011
elsif count = 177 then count <= 178; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 85, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 41, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 172, 8)),
6 => std_logic_vector(to_unsigned( 206, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 82, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 61, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 178 then count <= 179; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 37, 8)),
2 => std_logic_vector(to_unsigned( 4, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 41, 8)),
6 => std_logic_vector(to_unsigned( 83, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 66, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 179 then count <= 180; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 121, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 218, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 35, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 37, 8)),
10 => std_logic_vector(to_unsigned( 56, 8)),
11 => std_logic_vector(to_unsigned( 226, 8)),
12 => std_logic_vector(to_unsigned( 37, 8)),
13 => std_logic_vector(to_unsigned( 20, 8)),
14 => std_logic_vector(to_unsigned( 75, 8)),
15 => std_logic_vector(to_unsigned( 21, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 180 then count <= 181; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 254, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 2, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 242, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 232, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 215, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 213, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 181 then count <= 182; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 111, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 185, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 23, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 200, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 246, 8)),
16 => std_logic_vector(to_unsigned( 252, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 182 then count <= 183; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 5, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 21, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 225, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 166, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 189, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 205, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 183 then count <= 184; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 23, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 32, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 221, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 192, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 191, 8)),
16 => std_logic_vector(to_unsigned( 13, 8)),
17 => std_logic_vector(to_unsigned( 184, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 184 then count <= 185; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 24, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 108, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 41, 8)),
9 => std_logic_vector(to_unsigned( 31, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 24, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 104, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 185 then count <= 186; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 49, 8)),
4 => std_logic_vector(to_unsigned( 193, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 95, 8)),
14 => std_logic_vector(to_unsigned( 185, 8)),
15 => std_logic_vector(to_unsigned( 10, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 186 then count <= 187; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 6, 8)),
3 => std_logic_vector(to_unsigned( 21, 8)),
4 => std_logic_vector(to_unsigned( 247, 8)),
5 => std_logic_vector(to_unsigned( 133, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 168, 8)),
8 => std_logic_vector(to_unsigned( 233, 8)),
9 => std_logic_vector(to_unsigned( 184, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 187 then count <= 188; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 27, 8)),
2 => std_logic_vector(to_unsigned( 252, 8)),
3 => std_logic_vector(to_unsigned( 112, 8)),
4 => std_logic_vector(to_unsigned( 15, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 112, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 48, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 215, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 188 then count <= 189; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 49, 8)),
2 => std_logic_vector(to_unsigned( 202, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 245, 8)),
8 => std_logic_vector(to_unsigned( 91, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 57, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 70, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110010
elsif count = 189 then count <= 190; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 66, 8)),
2 => std_logic_vector(to_unsigned( 157, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 61, 8)),
6 => std_logic_vector(to_unsigned( 68, 8)),
7 => std_logic_vector(to_unsigned( 24, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 38, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 46, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 14, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 190 then count <= 191; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 169, 8)),
3 => std_logic_vector(to_unsigned( 21, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 158, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 169, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 185, 8)),
13 => std_logic_vector(to_unsigned( 228, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 0, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 191 then count <= 192; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 149, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 139, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 224, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 183, 8)),
14 => std_logic_vector(to_unsigned( 182, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 75, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 192 then count <= 193; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 200, 8)),
7 => std_logic_vector(to_unsigned( 254, 8)),
8 => std_logic_vector(to_unsigned( 2, 8)),
9 => std_logic_vector(to_unsigned( 206, 8)),
10 => std_logic_vector(to_unsigned( 180, 8)),
11 => std_logic_vector(to_unsigned( 254, 8)),
12 => std_logic_vector(to_unsigned( 40, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 243, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 241, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 183, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 193 then count <= 194; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 211, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 182, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 204, 8)),
9 => std_logic_vector(to_unsigned( 217, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 136, 8)),
12 => std_logic_vector(to_unsigned( 219, 8)),
13 => std_logic_vector(to_unsigned( 192, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 194 then count <= 195; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 47, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 103, 8)),
7 => std_logic_vector(to_unsigned( 133, 8)),
8 => std_logic_vector(to_unsigned( 20, 8)),
9 => std_logic_vector(to_unsigned( 5, 8)),
10 => std_logic_vector(to_unsigned( 15, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 217, 8)),
13 => std_logic_vector(to_unsigned( 24, 8)),
14 => std_logic_vector(to_unsigned( 146, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001101
elsif count = 195 then count <= 196; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 9, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 230, 8)),
10 => std_logic_vector(to_unsigned( 139, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 177, 8)),
15 => std_logic_vector(to_unsigned( 204, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 196 then count <= 197; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 62, 8)),
2 => std_logic_vector(to_unsigned( 192, 8)),
3 => std_logic_vector(to_unsigned( 73, 8)),
4 => std_logic_vector(to_unsigned( 165, 8)),
5 => std_logic_vector(to_unsigned( 20, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 130, 8)),
10 => std_logic_vector(to_unsigned( 214, 8)),
11 => std_logic_vector(to_unsigned( 36, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 9, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 134, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010011
elsif count = 197 then count <= 198; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 100, 8)),
4 => std_logic_vector(to_unsigned( 88, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 146, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 250, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 130, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 198 then count <= 199; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 45, 8)),
4 => std_logic_vector(to_unsigned( 14, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 249, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 95, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 183, 8)),
14 => std_logic_vector(to_unsigned( 205, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 184, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 199 then count <= 200; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 59, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 154, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 186, 8)),
13 => std_logic_vector(to_unsigned( 253, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 73, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 200 then count <= 201; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 18, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 13, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 62, 8)),
12 => std_logic_vector(to_unsigned( 227, 8)),
13 => std_logic_vector(to_unsigned( 15, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 23, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 201 then count <= 202; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 220, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 23, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 75, 8)),
11 => std_logic_vector(to_unsigned( 211, 8)),
12 => std_logic_vector(to_unsigned( 165, 8)),
13 => std_logic_vector(to_unsigned( 223, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 215, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 202 then count <= 203; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 176, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 59, 8)),
6 => std_logic_vector(to_unsigned( 197, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 195, 8)),
11 => std_logic_vector(to_unsigned( 78, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 255, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 203 then count <= 204; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 241, 8)),
2 => std_logic_vector(to_unsigned( 11, 8)),
3 => std_logic_vector(to_unsigned( 196, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 52, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 220, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 204 then count <= 205; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 5, 8)),
3 => std_logic_vector(to_unsigned( 98, 8)),
4 => std_logic_vector(to_unsigned( 45, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 148, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 42, 8)),
10 => std_logic_vector(to_unsigned( 236, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 16, 8)),
13 => std_logic_vector(to_unsigned( 181, 8)),
14 => std_logic_vector(to_unsigned( 50, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 49, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 205 then count <= 206; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 146, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 203, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 249, 8)),
8 => std_logic_vector(to_unsigned( 249, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 171, 8)),
15 => std_logic_vector(to_unsigned( 180, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 128, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 206 then count <= 207; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 16, 8)),
5 => std_logic_vector(to_unsigned( 8, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 34, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 204, 8)),
12 => std_logic_vector(to_unsigned( 37, 8)),
13 => std_logic_vector(to_unsigned( 200, 8)),
14 => std_logic_vector(to_unsigned( 67, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 108, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 50, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 207 then count <= 208; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 62, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 24, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 215, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 96, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 105, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 208 then count <= 209; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 101, 8)),
4 => std_logic_vector(to_unsigned( 228, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 244, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 135, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 68, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 238, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 209 then count <= 210; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 82, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 164, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 26, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 188, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 210 then count <= 211; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 55, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 147, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 156, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 211 then count <= 212; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 239, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 131, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 234, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 212 then count <= 213; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 57, 8)),
3 => std_logic_vector(to_unsigned( 55, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 249, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 20, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 82, 8)),
10 => std_logic_vector(to_unsigned( 124, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 223, 8)),
13 => std_logic_vector(to_unsigned( 55, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 5, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 213 then count <= 214; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 24, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 226, 8)),
6 => std_logic_vector(to_unsigned( 18, 8)),
7 => std_logic_vector(to_unsigned( 141, 8)),
8 => std_logic_vector(to_unsigned( 241, 8)),
9 => std_logic_vector(to_unsigned( 199, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 187, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 214 then count <= 215; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 49, 8)),
2 => std_logic_vector(to_unsigned( 200, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 52, 8)),
6 => std_logic_vector(to_unsigned( 197, 8)),
7 => std_logic_vector(to_unsigned( 38, 8)),
8 => std_logic_vector(to_unsigned( 127, 8)),
9 => std_logic_vector(to_unsigned( 145, 8)),
10 => std_logic_vector(to_unsigned( 48, 8)),
11 => std_logic_vector(to_unsigned( 76, 8)),
12 => std_logic_vector(to_unsigned( 235, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 248, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 61, 8)),
18 => std_logic_vector(to_unsigned( 219, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 215 then count <= 216; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 141, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 248, 8)),
5 => std_logic_vector(to_unsigned( 218, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 231, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 66, 8)),
14 => std_logic_vector(to_unsigned( 229, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 103, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 216 then count <= 217; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 203, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 39, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 30, 8)),
9 => std_logic_vector(to_unsigned( 199, 8)),
10 => std_logic_vector(to_unsigned( 1, 8)),
11 => std_logic_vector(to_unsigned( 193, 8)),
12 => std_logic_vector(to_unsigned( 71, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 66, 8)),
15 => std_logic_vector(to_unsigned( 74, 8)),
16 => std_logic_vector(to_unsigned( 52, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 39, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 217 then count <= 218; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 214, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 32, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 64, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 218 then count <= 219; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 153, 8)),
3 => std_logic_vector(to_unsigned( 208, 8)),
4 => std_logic_vector(to_unsigned( 89, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 189, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 254, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 151, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 219 then count <= 220; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 95, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 75, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 85, 8)),
6 => std_logic_vector(to_unsigned( 142, 8)),
7 => std_logic_vector(to_unsigned( 6, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 22, 8)),
11 => std_logic_vector(to_unsigned( 209, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 50, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 220 then count <= 221; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 0, 8)),
6 => std_logic_vector(to_unsigned( 87, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 238, 8)),
10 => std_logic_vector(to_unsigned( 59, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 13, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 168, 8)),
16 => std_logic_vector(to_unsigned( 108, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 221 then count <= 222; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 180, 8)),
6 => std_logic_vector(to_unsigned( 68, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 16, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 30, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 69, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 196, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 222 then count <= 223; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 120, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 251, 8)),
11 => std_logic_vector(to_unsigned( 246, 8)),
12 => std_logic_vector(to_unsigned( 157, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 239, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 213, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 223 then count <= 224; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 43, 8)),
2 => std_logic_vector(to_unsigned( 45, 8)),
3 => std_logic_vector(to_unsigned( 209, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 130, 8)),
10 => std_logic_vector(to_unsigned( 70, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 37, 8)),
15 => std_logic_vector(to_unsigned( 229, 8)),
16 => std_logic_vector(to_unsigned( 108, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 224 then count <= 225; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 236, 8)),
2 => std_logic_vector(to_unsigned( 94, 8)),
3 => std_logic_vector(to_unsigned( 79, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 197, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 34, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 131, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 210, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 11, 8)),
17 => std_logic_vector(to_unsigned( 188, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 225 then count <= 226; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 210, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 117, 8)),
5 => std_logic_vector(to_unsigned( 205, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 95, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 248, 8)),
14 => std_logic_vector(to_unsigned( 209, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 57, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 226 then count <= 227; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 168, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 201, 8)),
4 => std_logic_vector(to_unsigned( 41, 8)),
5 => std_logic_vector(to_unsigned( 46, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 216, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 6, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 32, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001010
elsif count = 227 then count <= 228; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 198, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 153, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 173, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 221, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 153, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 37, 8)),
14 => std_logic_vector(to_unsigned( 12, 8)),
15 => std_logic_vector(to_unsigned( 233, 8)),
16 => std_logic_vector(to_unsigned( 241, 8)),
17 => std_logic_vector(to_unsigned( 190, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 228 then count <= 229; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 139, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 199, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 220, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 135, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 195, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 199, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 229 then count <= 230; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 55, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 15, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 58, 8)),
9 => std_logic_vector(to_unsigned( 252, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 132, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 230 then count <= 231; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 49, 8)),
5 => std_logic_vector(to_unsigned( 29, 8)),
6 => std_logic_vector(to_unsigned( 50, 8)),
7 => std_logic_vector(to_unsigned( 218, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 84, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 10, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 136, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 231 then count <= 232; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 236, 8)),
3 => std_logic_vector(to_unsigned( 186, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 18, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 58, 8)),
9 => std_logic_vector(to_unsigned( 141, 8)),
10 => std_logic_vector(to_unsigned( 32, 8)),
11 => std_logic_vector(to_unsigned( 85, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 143, 8)),
16 => std_logic_vector(to_unsigned( 60, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 45, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 232 then count <= 233; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 219, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 77, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 172, 8)),
15 => std_logic_vector(to_unsigned( 45, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 57, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 233 then count <= 234; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 184, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 248, 8)),
10 => std_logic_vector(to_unsigned( 162, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 29, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 234 then count <= 235; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 204, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 54, 8)),
5 => std_logic_vector(to_unsigned( 245, 8)),
6 => std_logic_vector(to_unsigned( 202, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 60, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 100, 8)),
15 => std_logic_vector(to_unsigned( 61, 8)),
16 => std_logic_vector(to_unsigned( 51, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 64, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 235 then count <= 236; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 217, 8)),
2 => std_logic_vector(to_unsigned( 38, 8)),
3 => std_logic_vector(to_unsigned( 79, 8)),
4 => std_logic_vector(to_unsigned( 45, 8)),
5 => std_logic_vector(to_unsigned( 208, 8)),
6 => std_logic_vector(to_unsigned( 29, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 218, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 12, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 223, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 203, 8)),
18 => std_logic_vector(to_unsigned( 60, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 236 then count <= 237; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 155, 8)),
2 => std_logic_vector(to_unsigned( 200, 8)),
3 => std_logic_vector(to_unsigned( 19, 8)),
4 => std_logic_vector(to_unsigned( 106, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 184, 8)),
7 => std_logic_vector(to_unsigned( 11, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 230, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 173, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 219, 8)),
15 => std_logic_vector(to_unsigned( 128, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 237 then count <= 238; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 68, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 113, 8)),
4 => std_logic_vector(to_unsigned( 224, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 216, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 179, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 182, 8)),
13 => std_logic_vector(to_unsigned( 221, 8)),
14 => std_logic_vector(to_unsigned( 229, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 193, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 238 then count <= 239; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 14, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 152, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 239 then count <= 240; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 15, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 230, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 22, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 20, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 240 then count <= 241; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 40, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 29, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 30, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 181, 8)),
12 => std_logic_vector(to_unsigned( 36, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 79, 8)),
17 => std_logic_vector(to_unsigned( 39, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 241 then count <= 242; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 9, 8)),
2 => std_logic_vector(to_unsigned( 57, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 23, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 242 then count <= 243; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 37, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 230, 8)),
5 => std_logic_vector(to_unsigned( 230, 8)),
6 => std_logic_vector(to_unsigned( 212, 8)),
7 => std_logic_vector(to_unsigned( 27, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 16, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 243 then count <= 244; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 18, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 73, 8)),
7 => std_logic_vector(to_unsigned( 66, 8)),
8 => std_logic_vector(to_unsigned( 55, 8)),
9 => std_logic_vector(to_unsigned( 156, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 15, 8)),
12 => std_logic_vector(to_unsigned( 189, 8)),
13 => std_logic_vector(to_unsigned( 151, 8)),
14 => std_logic_vector(to_unsigned( 80, 8)),
15 => std_logic_vector(to_unsigned( 40, 8)),
16 => std_logic_vector(to_unsigned( 97, 8)),
17 => std_logic_vector(to_unsigned( 40, 8)),
18 => std_logic_vector(to_unsigned( 63, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 244 then count <= 245; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 237, 8)),
2 => std_logic_vector(to_unsigned( 155, 8)),
3 => std_logic_vector(to_unsigned( 59, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 228, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 212, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 185, 8)),
17 => std_logic_vector(to_unsigned( 218, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 245 then count <= 246; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 49, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 220, 8)),
5 => std_logic_vector(to_unsigned( 112, 8)),
6 => std_logic_vector(to_unsigned( 231, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 188, 8)),
10 => std_logic_vector(to_unsigned( 12, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 138, 8)),
13 => std_logic_vector(to_unsigned( 235, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 246 then count <= 247; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 150, 8)),
12 => std_logic_vector(to_unsigned( 154, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 247 then count <= 248; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 155, 8)),
2 => std_logic_vector(to_unsigned( 142, 8)),
3 => std_logic_vector(to_unsigned( 221, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 250, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 214, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 188, 8)),
12 => std_logic_vector(to_unsigned( 109, 8)),
13 => std_logic_vector(to_unsigned( 195, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 56, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 248 then count <= 249; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 223, 8)),
2 => std_logic_vector(to_unsigned( 61, 8)),
3 => std_logic_vector(to_unsigned( 63, 8)),
4 => std_logic_vector(to_unsigned( 228, 8)),
5 => std_logic_vector(to_unsigned( 198, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 237, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 216, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 16, 8)),
13 => std_logic_vector(to_unsigned( 185, 8)),
14 => std_logic_vector(to_unsigned( 135, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 210, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 249 then count <= 250; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 233, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 35, 8)),
4 => std_logic_vector(to_unsigned( 89, 8)),
5 => std_logic_vector(to_unsigned( 9, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 101, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 119, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 250 then count <= 251; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 195, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 106, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 148, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 17, 8)),
16 => std_logic_vector(to_unsigned( 25, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 251 then count <= 252; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 25, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 68, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 68, 8)),
11 => std_logic_vector(to_unsigned( 55, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 82, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 63, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 252 then count <= 253; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 215, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 255, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 50, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 253 then count <= 254; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 24, 8)),
3 => std_logic_vector(to_unsigned( 248, 8)),
4 => std_logic_vector(to_unsigned( 166, 8)),
5 => std_logic_vector(to_unsigned( 192, 8)),
6 => std_logic_vector(to_unsigned( 6, 8)),
7 => std_logic_vector(to_unsigned( 189, 8)),
8 => std_logic_vector(to_unsigned( 9, 8)),
9 => std_logic_vector(to_unsigned( 13, 8)),
10 => std_logic_vector(to_unsigned( 35, 8)),
11 => std_logic_vector(to_unsigned( 205, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 232, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 237, 8)),
16 => std_logic_vector(to_unsigned( 43, 8)),
17 => std_logic_vector(to_unsigned( 196, 8)),
18 => std_logic_vector(to_unsigned( 44, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 254 then count <= 255; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 253, 8)),
2 => std_logic_vector(to_unsigned( 64, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 202, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 139, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 97, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 255 then count <= 256; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 241, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 85, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 221, 8)),
8 => std_logic_vector(to_unsigned( 42, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 251, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 256 then count <= 257; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 198, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 146, 8)),
6 => std_logic_vector(to_unsigned( 175, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 13, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 222, 8)),
13 => std_logic_vector(to_unsigned( 87, 8)),
14 => std_logic_vector(to_unsigned( 185, 8)),
15 => std_logic_vector(to_unsigned( 80, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00100111
elsif count = 257 then count <= 258; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 239, 8)),
5 => std_logic_vector(to_unsigned( 193, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 180, 8)),
8 => std_logic_vector(to_unsigned( 211, 8)),
9 => std_logic_vector(to_unsigned( 0, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 223, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 258 then count <= 259; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 94, 8)),
3 => std_logic_vector(to_unsigned( 195, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 59, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 46, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 248, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 56, 8)),
15 => std_logic_vector(to_unsigned( 214, 8)),
16 => std_logic_vector(to_unsigned( 51, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 259 then count <= 260; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 157, 8)),
3 => std_logic_vector(to_unsigned( 74, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 89, 8)),
8 => std_logic_vector(to_unsigned( 211, 8)),
9 => std_logic_vector(to_unsigned( 241, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001011
elsif count = 260 then count <= 261; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 182, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 201, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 261 then count <= 262; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 68, 8)),
2 => std_logic_vector(to_unsigned( 211, 8)),
3 => std_logic_vector(to_unsigned( 226, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 245, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 15, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 136, 8)),
14 => std_logic_vector(to_unsigned( 135, 8)),
15 => std_logic_vector(to_unsigned( 233, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 262 then count <= 263; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 110, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 244, 8)),
8 => std_logic_vector(to_unsigned( 60, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 113, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 263 then count <= 264; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 118, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 8, 8)),
8 => std_logic_vector(to_unsigned( 251, 8)),
9 => std_logic_vector(to_unsigned( 89, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 23, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 28, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 264 then count <= 265; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 229, 8)),
4 => std_logic_vector(to_unsigned( 14, 8)),
5 => std_logic_vector(to_unsigned( 112, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 20, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 47, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 56, 8)),
16 => std_logic_vector(to_unsigned( 95, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 265 then count <= 266; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 29, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 98, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 19, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 52, 8)),
8 => std_logic_vector(to_unsigned( 249, 8)),
9 => std_logic_vector(to_unsigned( 33, 8)),
10 => std_logic_vector(to_unsigned( 217, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 228, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 86, 8)),
16 => std_logic_vector(to_unsigned( 210, 8)),
17 => std_logic_vector(to_unsigned( 56, 8)),
18 => std_logic_vector(to_unsigned( 197, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 266 then count <= 267; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 116, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 125, 8)),
7 => std_logic_vector(to_unsigned( 83, 8)),
8 => std_logic_vector(to_unsigned( 155, 8)),
9 => std_logic_vector(to_unsigned( 134, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 215, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 39, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 187, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 133, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 267 then count <= 268; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 51, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 208, 8)),
14 => std_logic_vector(to_unsigned( 41, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 268 then count <= 269; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 165, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 244, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 176, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 138, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 269 then count <= 270; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 19, 8)),
3 => std_logic_vector(to_unsigned( 109, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 33, 8)),
6 => std_logic_vector(to_unsigned( 59, 8)),
7 => std_logic_vector(to_unsigned( 67, 8)),
8 => std_logic_vector(to_unsigned( 25, 8)),
9 => std_logic_vector(to_unsigned( 156, 8)),
10 => std_logic_vector(to_unsigned( 68, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 254, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 270 then count <= 271; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 81, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 125, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 214, 8)),
10 => std_logic_vector(to_unsigned( 248, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 252, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 271 then count <= 272; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 231, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 272 then count <= 273; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 91, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 137, 8)),
7 => std_logic_vector(to_unsigned( 4, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 71, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 212, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 273 then count <= 274; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 15, 8)),
5 => std_logic_vector(to_unsigned( 251, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 23, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 34, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 102, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 274 then count <= 275; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 144, 8)),
3 => std_logic_vector(to_unsigned( 190, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 189, 8)),
6 => std_logic_vector(to_unsigned( 248, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 58, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 100, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 275 then count <= 276; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 224, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 91, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 141, 8)),
10 => std_logic_vector(to_unsigned( 216, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 213, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 46, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 276 then count <= 277; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 238, 8)),
2 => std_logic_vector(to_unsigned( 238, 8)),
3 => std_logic_vector(to_unsigned( 222, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 219, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 223, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 219, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 277 then count <= 278; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 31, 8)),
2 => std_logic_vector(to_unsigned( 241, 8)),
3 => std_logic_vector(to_unsigned( 211, 8)),
4 => std_logic_vector(to_unsigned( 240, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 132, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 216, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011000
elsif count = 278 then count <= 279; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 129, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 28, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 80, 8)),
10 => std_logic_vector(to_unsigned( 234, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 225, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 128, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 213, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 279 then count <= 280; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 10, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 54, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 178, 8)),
15 => std_logic_vector(to_unsigned( 32, 8)),
16 => std_logic_vector(to_unsigned( 103, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 280 then count <= 281; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 94, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 182, 8)),
11 => std_logic_vector(to_unsigned( 83, 8)),
12 => std_logic_vector(to_unsigned( 193, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 214, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 281 then count <= 282; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 196, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 203, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 149, 8)),
6 => std_logic_vector(to_unsigned( 127, 8)),
7 => std_logic_vector(to_unsigned( 248, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 229, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 145, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 282 then count <= 283; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 240, 8)),
6 => std_logic_vector(to_unsigned( 231, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 137, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 105, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 56, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 283 then count <= 284; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 155, 8)),
2 => std_logic_vector(to_unsigned( 131, 8)),
3 => std_logic_vector(to_unsigned( 234, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 20, 8)),
12 => std_logic_vector(to_unsigned( 58, 8)),
13 => std_logic_vector(to_unsigned( 133, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 25, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 284 then count <= 285; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 158, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 105, 8)),
5 => std_logic_vector(to_unsigned( 9, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 213, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 228, 8)),
10 => std_logic_vector(to_unsigned( 142, 8)),
11 => std_logic_vector(to_unsigned( 19, 8)),
12 => std_logic_vector(to_unsigned( 154, 8)),
13 => std_logic_vector(to_unsigned( 201, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 285 then count <= 286; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 28, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 34, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 243, 8)),
7 => std_logic_vector(to_unsigned( 53, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 54, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 128, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 286 then count <= 287; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 26, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 163, 8)),
6 => std_logic_vector(to_unsigned( 231, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 193, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 199, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 30, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 287 then count <= 288; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 194, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 155, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 186, 8)),
9 => std_logic_vector(to_unsigned( 11, 8)),
10 => std_logic_vector(to_unsigned( 190, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 102, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 288 then count <= 289; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 127, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 78, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 224, 8)),
13 => std_logic_vector(to_unsigned( 186, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 173, 8)),
16 => std_logic_vector(to_unsigned( 230, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 289 then count <= 290; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 235, 8)),
2 => std_logic_vector(to_unsigned( 234, 8)),
3 => std_logic_vector(to_unsigned( 19, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 68, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 90, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 211, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 179, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 290 then count <= 291; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 191, 8)),
3 => std_logic_vector(to_unsigned( 150, 8)),
4 => std_logic_vector(to_unsigned( 10, 8)),
5 => std_logic_vector(to_unsigned( 170, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 21, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 228, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 33, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 291 then count <= 292; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 37, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 192, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 175, 8)),
11 => std_logic_vector(to_unsigned( 16, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 250, 8)),
14 => std_logic_vector(to_unsigned( 16, 8)),
15 => std_logic_vector(to_unsigned( 136, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 73, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 292 then count <= 293; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 190, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 21, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 249, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 45, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 170, 8)),
14 => std_logic_vector(to_unsigned( 41, 8)),
15 => std_logic_vector(to_unsigned( 172, 8)),
16 => std_logic_vector(to_unsigned( 43, 8)),
17 => std_logic_vector(to_unsigned( 210, 8)),
18 => std_logic_vector(to_unsigned( 41, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 293 then count <= 294; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 118, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 11, 8)),
5 => std_logic_vector(to_unsigned( 28, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 135, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 163, 8)),
12 => std_logic_vector(to_unsigned( 46, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 45, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100010
elsif count = 294 then count <= 295; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 58, 8)),
2 => std_logic_vector(to_unsigned( 9, 8)),
3 => std_logic_vector(to_unsigned( 237, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 255, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 237, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 30, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 92, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 295 then count <= 296; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 5, 8)),
11 => std_logic_vector(to_unsigned( 204, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 226, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 296 then count <= 297; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 198, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 241, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 28, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 47, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 297 then count <= 298; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 75, 8)),
5 => std_logic_vector(to_unsigned( 182, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 181, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 159, 8)),
12 => std_logic_vector(to_unsigned( 242, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 298 then count <= 299; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 165, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 17, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 189, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 244, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 196, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 199, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 299 then count <= 300; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 27, 8)),
3 => std_logic_vector(to_unsigned( 16, 8)),
4 => std_logic_vector(to_unsigned( 240, 8)),
5 => std_logic_vector(to_unsigned( 46, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 172, 8)),
16 => std_logic_vector(to_unsigned( 49, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 300 then count <= 301; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 230, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 301 then count <= 302; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 71, 8)),
3 => std_logic_vector(to_unsigned( 251, 8)),
4 => std_logic_vector(to_unsigned( 38, 8)),
5 => std_logic_vector(to_unsigned( 115, 8)),
6 => std_logic_vector(to_unsigned( 4, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 216, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 31, 8)),
13 => std_logic_vector(to_unsigned( 39, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 103, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 53, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110101
elsif count = 302 then count <= 303; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 81, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 241, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 63, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 207, 8)),
14 => std_logic_vector(to_unsigned( 28, 8)),
15 => std_logic_vector(to_unsigned( 46, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 303 then count <= 304; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 220, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 21, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 188, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 26, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 55, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110110
elsif count = 304 then count <= 305; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 78, 8)),
5 => std_logic_vector(to_unsigned( 55, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 26, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 27, 8)),
11 => std_logic_vector(to_unsigned( 107, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 40, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 32, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 305 then count <= 306; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 185, 8)),
2 => std_logic_vector(to_unsigned( 242, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 240, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 170, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 228, 8)),
17 => std_logic_vector(to_unsigned( 184, 8)),
18 => std_logic_vector(to_unsigned( 210, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 306 then count <= 307; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 130, 8)),
2 => std_logic_vector(to_unsigned( 9, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 123, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 88, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 196, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 71, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 307 then count <= 308; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 8, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 224, 8)),
5 => std_logic_vector(to_unsigned( 82, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 137, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 6, 8)),
14 => std_logic_vector(to_unsigned( 250, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 308 then count <= 309; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 56, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 32, 8)),
7 => std_logic_vector(to_unsigned( 21, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 107, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 152, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 59, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 309 then count <= 310; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 176, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 90, 8)),
5 => std_logic_vector(to_unsigned( 117, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 41, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 85, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 173, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 310 then count <= 311; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 27, 8)),
6 => std_logic_vector(to_unsigned( 53, 8)),
7 => std_logic_vector(to_unsigned( 42, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 86, 8)),
12 => std_logic_vector(to_unsigned( 36, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 311 then count <= 312; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 18, 8)),
3 => std_logic_vector(to_unsigned( 15, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 144, 8)),
9 => std_logic_vector(to_unsigned( 45, 8)),
10 => std_logic_vector(to_unsigned( 197, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 27, 8)),
13 => std_logic_vector(to_unsigned( 18, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 312 then count <= 313; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 64, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 248, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 28, 8)),
10 => std_logic_vector(to_unsigned( 108, 8)),
11 => std_logic_vector(to_unsigned( 54, 8)),
12 => std_logic_vector(to_unsigned( 39, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 77, 8)),
15 => std_logic_vector(to_unsigned( 236, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00010111
elsif count = 313 then count <= 314; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 200, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 229, 8)),
8 => std_logic_vector(to_unsigned( 49, 8)),
9 => std_logic_vector(to_unsigned( 206, 8)),
10 => std_logic_vector(to_unsigned( 79, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 60, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 314 then count <= 315; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 60, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 211, 8)),
6 => std_logic_vector(to_unsigned( 68, 8)),
7 => std_logic_vector(to_unsigned( 202, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 240, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 191, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 237, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 172, 8)),
16 => std_logic_vector(to_unsigned( 18, 8)),
17 => std_logic_vector(to_unsigned( 202, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 315 then count <= 316; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 198, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 232, 8)),
4 => std_logic_vector(to_unsigned( 71, 8)),
5 => std_logic_vector(to_unsigned( 44, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 207, 8)),
8 => std_logic_vector(to_unsigned( 40, 8)),
9 => std_logic_vector(to_unsigned( 19, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 249, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 316 then count <= 317; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 216, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 213, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 219, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 24, 8)),
14 => std_logic_vector(to_unsigned( 254, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 14, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 317 then count <= 318; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 47, 8)),
2 => std_logic_vector(to_unsigned( 143, 8)),
3 => std_logic_vector(to_unsigned( 20, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 195, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 15, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 23, 8)),
14 => std_logic_vector(to_unsigned( 41, 8)),
15 => std_logic_vector(to_unsigned( 31, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 37, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 318 then count <= 319; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 235, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 156, 8)),
7 => std_logic_vector(to_unsigned( 60, 8)),
8 => std_logic_vector(to_unsigned( 109, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 180, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 214, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 319 then count <= 320; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 176, 8)),
3 => std_logic_vector(to_unsigned( 253, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 155, 8)),
14 => std_logic_vector(to_unsigned( 236, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 320 then count <= 321; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 248, 8)),
2 => std_logic_vector(to_unsigned( 54, 8)),
3 => std_logic_vector(to_unsigned( 120, 8)),
4 => std_logic_vector(to_unsigned( 185, 8)),
5 => std_logic_vector(to_unsigned( 184, 8)),
6 => std_logic_vector(to_unsigned( 216, 8)),
7 => std_logic_vector(to_unsigned( 84, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 69, 8)),
12 => std_logic_vector(to_unsigned( 110, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 35, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 321 then count <= 322; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 169, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 132, 8)),
8 => std_logic_vector(to_unsigned( 82, 8)),
9 => std_logic_vector(to_unsigned( 28, 8)),
10 => std_logic_vector(to_unsigned( 36, 8)),
11 => std_logic_vector(to_unsigned( 36, 8)),
12 => std_logic_vector(to_unsigned( 182, 8)),
13 => std_logic_vector(to_unsigned( 196, 8)),
14 => std_logic_vector(to_unsigned( 128, 8)),
15 => std_logic_vector(to_unsigned( 212, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 322 then count <= 323; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 243, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 208, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110010
elsif count = 323 then count <= 324; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 248, 8)),
3 => std_logic_vector(to_unsigned( 108, 8)),
4 => std_logic_vector(to_unsigned( 79, 8)),
5 => std_logic_vector(to_unsigned( 86, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 77, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 324 then count <= 325; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 72, 8)),
2 => std_logic_vector(to_unsigned( 21, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 61, 8)),
5 => std_logic_vector(to_unsigned( 25, 8)),
6 => std_logic_vector(to_unsigned( 15, 8)),
7 => std_logic_vector(to_unsigned( 39, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 70, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 59, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101010
elsif count = 325 then count <= 326; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 122, 8)),
6 => std_logic_vector(to_unsigned( 207, 8)),
7 => std_logic_vector(to_unsigned( 60, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 74, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 201, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 133, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 326 then count <= 327; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 200, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 157, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 10, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 327 then count <= 328; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 182, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 186, 8)),
9 => std_logic_vector(to_unsigned( 241, 8)),
10 => std_logic_vector(to_unsigned( 76, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 203, 8)),
13 => std_logic_vector(to_unsigned( 225, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 54, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 328 then count <= 329; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 141, 8)),
3 => std_logic_vector(to_unsigned( 224, 8)),
4 => std_logic_vector(to_unsigned( 173, 8)),
5 => std_logic_vector(to_unsigned( 216, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 216, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 46, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 329 then count <= 330; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 209, 8)),
4 => std_logic_vector(to_unsigned( 209, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 210, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 219, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 330 then count <= 331; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 20, 8)),
2 => std_logic_vector(to_unsigned( 136, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 166, 8)),
8 => std_logic_vector(to_unsigned( 185, 8)),
9 => std_logic_vector(to_unsigned( 224, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 216, 8)),
14 => std_logic_vector(to_unsigned( 144, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100010
elsif count = 331 then count <= 332; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 70, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 12, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 87, 8)),
11 => std_logic_vector(to_unsigned( 252, 8)),
12 => std_logic_vector(to_unsigned( 30, 8)),
13 => std_logic_vector(to_unsigned( 233, 8)),
14 => std_logic_vector(to_unsigned( 186, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 54, 8)),
17 => std_logic_vector(to_unsigned( 47, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 332 then count <= 333; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 251, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 227, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 164, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 41, 8)),
8 => std_logic_vector(to_unsigned( 193, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 131, 8)),
13 => std_logic_vector(to_unsigned( 152, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 333 then count <= 334; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 71, 8)),
3 => std_logic_vector(to_unsigned( 5, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 29, 8)),
6 => std_logic_vector(to_unsigned( 134, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 75, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 59, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 334 then count <= 335; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 67, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 194, 8)),
16 => std_logic_vector(to_unsigned( 230, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 335 then count <= 336; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 41, 8)),
4 => std_logic_vector(to_unsigned( 73, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 24, 8)),
7 => std_logic_vector(to_unsigned( 221, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 6, 8)),
12 => std_logic_vector(to_unsigned( 28, 8)),
13 => std_logic_vector(to_unsigned( 217, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 336 then count <= 337; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 62, 8)),
3 => std_logic_vector(to_unsigned( 181, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 183, 8)),
6 => std_logic_vector(to_unsigned( 199, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 68, 8)),
11 => std_logic_vector(to_unsigned( 210, 8)),
12 => std_logic_vector(to_unsigned( 234, 8)),
13 => std_logic_vector(to_unsigned( 208, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 337 then count <= 338; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 227, 8)),
2 => std_logic_vector(to_unsigned( 195, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 209, 8)),
9 => std_logic_vector(to_unsigned( 248, 8)),
10 => std_logic_vector(to_unsigned( 55, 8)),
11 => std_logic_vector(to_unsigned( 120, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 223, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 338 then count <= 339; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 192, 8)),
3 => std_logic_vector(to_unsigned( 207, 8)),
4 => std_logic_vector(to_unsigned( 173, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 0, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 226, 8)),
13 => std_logic_vector(to_unsigned( 13, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 240, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 339 then count <= 340; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 67, 8)),
3 => std_logic_vector(to_unsigned( 100, 8)),
4 => std_logic_vector(to_unsigned( 55, 8)),
5 => std_logic_vector(to_unsigned( 238, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 119, 8)),
10 => std_logic_vector(to_unsigned( 36, 8)),
11 => std_logic_vector(to_unsigned( 255, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 62, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 63, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 340 then count <= 341; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 252, 8)),
2 => std_logic_vector(to_unsigned( 198, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 118, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 33, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 208, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 180, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 341 then count <= 342; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 108, 8)),
5 => std_logic_vector(to_unsigned( 72, 8)),
6 => std_logic_vector(to_unsigned( 74, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 22, 8)),
9 => std_logic_vector(to_unsigned( 4, 8)),
10 => std_logic_vector(to_unsigned( 244, 8)),
11 => std_logic_vector(to_unsigned( 70, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 13, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 342 then count <= 343; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 75, 8)),
9 => std_logic_vector(to_unsigned( 11, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 3, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 222, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 343 then count <= 344; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 75, 8)),
2 => std_logic_vector(to_unsigned( 212, 8)),
3 => std_logic_vector(to_unsigned( 12, 8)),
4 => std_logic_vector(to_unsigned( 244, 8)),
5 => std_logic_vector(to_unsigned( 53, 8)),
6 => std_logic_vector(to_unsigned( 190, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 70, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 6, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 57, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 190, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 344 then count <= 345; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 217, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 234, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 225, 8)),
15 => std_logic_vector(to_unsigned( 51, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 345 then count <= 346; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 180, 8)),
2 => std_logic_vector(to_unsigned( 216, 8)),
3 => std_logic_vector(to_unsigned( 16, 8)),
4 => std_logic_vector(to_unsigned( 28, 8)),
5 => std_logic_vector(to_unsigned( 243, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 207, 8)),
12 => std_logic_vector(to_unsigned( 217, 8)),
13 => std_logic_vector(to_unsigned( 195, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 255, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 346 then count <= 347; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 245, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 177, 8)),
5 => std_logic_vector(to_unsigned( 248, 8)),
6 => std_logic_vector(to_unsigned( 197, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 155, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 228, 8)),
14 => std_logic_vector(to_unsigned( 12, 8)),
15 => std_logic_vector(to_unsigned( 152, 8)),
16 => std_logic_vector(to_unsigned( 126, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 347 then count <= 348; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 203, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 170, 8)),
5 => std_logic_vector(to_unsigned( 50, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 150, 8)),
8 => std_logic_vector(to_unsigned( 235, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 249, 8)),
13 => std_logic_vector(to_unsigned( 44, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 38, 8)),
16 => std_logic_vector(to_unsigned( 244, 8)),
17 => std_logic_vector(to_unsigned( 39, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 348 then count <= 349; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 91, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 76, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 105, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 43, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 60, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 349 then count <= 350; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 28, 8)),
3 => std_logic_vector(to_unsigned( 197, 8)),
4 => std_logic_vector(to_unsigned( 63, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 78, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 13, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 81, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 8, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 33, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 45, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 350 then count <= 351; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 235, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 0, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 34, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 185, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110010
elsif count = 351 then count <= 352; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 59, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 24, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 24, 8)),
7 => std_logic_vector(to_unsigned( 209, 8)),
8 => std_logic_vector(to_unsigned( 207, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 23, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 28, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 244, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 352 then count <= 353; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 57, 8)),
3 => std_logic_vector(to_unsigned( 86, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 212, 8)),
9 => std_logic_vector(to_unsigned( 232, 8)),
10 => std_logic_vector(to_unsigned( 142, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 353 then count <= 354; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 11, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 19, 8)),
4 => std_logic_vector(to_unsigned( 78, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 1, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 201, 8)),
13 => std_logic_vector(to_unsigned( 0, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 23, 8)),
16 => std_logic_vector(to_unsigned( 74, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 354 then count <= 355; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 32, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 13, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 81, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 182, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 355 then count <= 356; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 254, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 93, 8)),
6 => std_logic_vector(to_unsigned( 218, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 166, 8)),
9 => std_logic_vector(to_unsigned( 7, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 61, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 185, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 356 then count <= 357; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 19, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 83, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 222, 8)),
14 => std_logic_vector(to_unsigned( 62, 8)),
15 => std_logic_vector(to_unsigned( 193, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 357 then count <= 358; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 158, 8)),
2 => std_logic_vector(to_unsigned( 130, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 199, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 214, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 358 then count <= 359; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 90, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 148, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 238, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 251, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 131, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 359 then count <= 360; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 59, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 116, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 82, 8)),
9 => std_logic_vector(to_unsigned( 24, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 27, 8)),
16 => std_logic_vector(to_unsigned( 205, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101110
elsif count = 360 then count <= 361; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 39, 8)),
2 => std_logic_vector(to_unsigned( 131, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 33, 8)),
7 => std_logic_vector(to_unsigned( 1, 8)),
8 => std_logic_vector(to_unsigned( 14, 8)),
9 => std_logic_vector(to_unsigned( 96, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 59, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 361 then count <= 362; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 21, 8)),
3 => std_logic_vector(to_unsigned( 32, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 107, 8)),
9 => std_logic_vector(to_unsigned( 201, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 188, 8)),
13 => std_logic_vector(to_unsigned( 43, 8)),
14 => std_logic_vector(to_unsigned( 140, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 49, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 362 then count <= 363; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 45, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 222, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 77, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 38, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 195, 8)),
15 => std_logic_vector(to_unsigned( 25, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 46, 8)),
18 => std_logic_vector(to_unsigned( 64, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010011
elsif count = 363 then count <= 364; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 45, 8)),
4 => std_logic_vector(to_unsigned( 203, 8)),
5 => std_logic_vector(to_unsigned( 14, 8)),
6 => std_logic_vector(to_unsigned( 74, 8)),
7 => std_logic_vector(to_unsigned( 5, 8)),
8 => std_logic_vector(to_unsigned( 4, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 73, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110101
elsif count = 364 then count <= 365; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 12, 8)),
5 => std_logic_vector(to_unsigned( 33, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 167, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 151, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 4, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 365 then count <= 366; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 72, 8)),
2 => std_logic_vector(to_unsigned( 72, 8)),
3 => std_logic_vector(to_unsigned( 68, 8)),
4 => std_logic_vector(to_unsigned( 223, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 103, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 52, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 107, 8)),
11 => std_logic_vector(to_unsigned( 44, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 90, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 366 then count <= 367; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 1, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 80, 8)),
4 => std_logic_vector(to_unsigned( 112, 8)),
5 => std_logic_vector(to_unsigned( 117, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 77, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 196, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 23, 8)),
16 => std_logic_vector(to_unsigned( 238, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 367 then count <= 368; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 172, 8)),
6 => std_logic_vector(to_unsigned( 185, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 70, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 368 then count <= 369; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 25, 8)),
3 => std_logic_vector(to_unsigned( 203, 8)),
4 => std_logic_vector(to_unsigned( 0, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 76, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 59, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101100
elsif count = 369 then count <= 370; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 236, 8)),
7 => std_logic_vector(to_unsigned( 183, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 108, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 370 then count <= 371; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 254, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 2, 8)),
5 => std_logic_vector(to_unsigned( 243, 8)),
6 => std_logic_vector(to_unsigned( 212, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 24, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 2, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 32, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111010
elsif count = 371 then count <= 372; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 238, 8)),
5 => std_logic_vector(to_unsigned( 232, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 200, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 41, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 193, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 372 then count <= 373; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 223, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 180, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 182, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 373 then count <= 374; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 147, 8)),
2 => std_logic_vector(to_unsigned( 236, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 164, 8)),
6 => std_logic_vector(to_unsigned( 235, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 188, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 32, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 374 then count <= 375; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 235, 8)),
2 => std_logic_vector(to_unsigned( 240, 8)),
3 => std_logic_vector(to_unsigned( 196, 8)),
4 => std_logic_vector(to_unsigned( 173, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 214, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 241, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 28, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 241, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 375 then count <= 376; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 91, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 227, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 93, 8)),
9 => std_logic_vector(to_unsigned( 184, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 66, 8)),
12 => std_logic_vector(to_unsigned( 227, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 224, 8)),
16 => std_logic_vector(to_unsigned( 75, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 376 then count <= 377; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 76, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 89, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 377 then count <= 378; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 220, 8)),
3 => std_logic_vector(to_unsigned( 20, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 78, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 11, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 378 then count <= 379; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 188, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 185, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 20, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 20, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 135, 8)),
15 => std_logic_vector(to_unsigned( 250, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 379 then count <= 380; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 62, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 220, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 162, 8)),
11 => std_logic_vector(to_unsigned( 181, 8)),
12 => std_logic_vector(to_unsigned( 185, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 75, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 380 then count <= 381; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 101, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 41, 8)),
8 => std_logic_vector(to_unsigned( 159, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 227, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 192, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 381 then count <= 382; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 47, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 208, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 198, 8)),
7 => std_logic_vector(to_unsigned( 2, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 215, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 56, 8)),
15 => std_logic_vector(to_unsigned( 155, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 382 then count <= 383; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 34, 8)),
4 => std_logic_vector(to_unsigned( 92, 8)),
5 => std_logic_vector(to_unsigned( 205, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 43, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 16, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 54, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 383 then count <= 384; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 242, 8)),
5 => std_logic_vector(to_unsigned( 36, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 18, 8)),
11 => std_logic_vector(to_unsigned( 27, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 52, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 384 then count <= 385; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 221, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 215, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 248, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 165, 8)),
11 => std_logic_vector(to_unsigned( 250, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 240, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 11, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 385 then count <= 386; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 180, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 18, 8)),
5 => std_logic_vector(to_unsigned( 122, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 18, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 29, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 211, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 386 then count <= 387; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 89, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 215, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 250, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 39, 8)),
13 => std_logic_vector(to_unsigned( 221, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 387 then count <= 388; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 78, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 182, 8)),
10 => std_logic_vector(to_unsigned( 177, 8)),
11 => std_logic_vector(to_unsigned( 254, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 207, 8)),
14 => std_logic_vector(to_unsigned( 216, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 388 then count <= 389; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 236, 8)),
2 => std_logic_vector(to_unsigned( 5, 8)),
3 => std_logic_vector(to_unsigned( 12, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 142, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 66, 8)),
9 => std_logic_vector(to_unsigned( 86, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 29, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 80, 8)),
16 => std_logic_vector(to_unsigned( 24, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 40, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 389 then count <= 390; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 241, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 253, 8)),
7 => std_logic_vector(to_unsigned( 22, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 33, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 51, 8)),
14 => std_logic_vector(to_unsigned( 220, 8)),
15 => std_logic_vector(to_unsigned( 239, 8)),
16 => std_logic_vector(to_unsigned( 17, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 390 then count <= 391; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 199, 8)),
2 => std_logic_vector(to_unsigned( 31, 8)),
3 => std_logic_vector(to_unsigned( 153, 8)),
4 => std_logic_vector(to_unsigned( 108, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 136, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 58, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 391 then count <= 392; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 19, 8)),
2 => std_logic_vector(to_unsigned( 196, 8)),
3 => std_logic_vector(to_unsigned( 63, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 198, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 163, 8)),
11 => std_logic_vector(to_unsigned( 72, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 20, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 392 then count <= 393; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 14, 8)),
2 => std_logic_vector(to_unsigned( 130, 8)),
3 => std_logic_vector(to_unsigned( 16, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 3, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 147, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 41, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 178, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 393 then count <= 394; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 215, 8)),
5 => std_logic_vector(to_unsigned( 103, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 209, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 394 then count <= 395; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 30, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 22, 8)),
5 => std_logic_vector(to_unsigned( 93, 8)),
6 => std_logic_vector(to_unsigned( 66, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 29, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 12, 8)),
13 => std_logic_vector(to_unsigned( 236, 8)),
14 => std_logic_vector(to_unsigned( 12, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110110
elsif count = 395 then count <= 396; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 42, 8)),
2 => std_logic_vector(to_unsigned( 239, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 27, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 209, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 240, 8)),
10 => std_logic_vector(to_unsigned( 212, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 96, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100100
elsif count = 396 then count <= 397; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 151, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 112, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 183, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 255, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 1, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010111
elsif count = 397 then count <= 398; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 172, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 189, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 141, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 213, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 182, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 398 then count <= 399; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 241, 8)),
4 => std_logic_vector(to_unsigned( 73, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 185, 8)),
7 => std_logic_vector(to_unsigned( 11, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 74, 8)),
15 => std_logic_vector(to_unsigned( 88, 8)),
16 => std_logic_vector(to_unsigned( 168, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110101
elsif count = 399 then count <= 400; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 250, 8)),
2 => std_logic_vector(to_unsigned( 197, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 21, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 49, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 18, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 400 then count <= 401; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 33, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 91, 8)),
6 => std_logic_vector(to_unsigned( 242, 8)),
7 => std_logic_vector(to_unsigned( 108, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 131, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 190, 8)),
14 => std_logic_vector(to_unsigned( 34, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 32, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 54, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 401 then count <= 402; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 232, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 241, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 22, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 59, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 85, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 173, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 402 then count <= 403; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 247, 8)),
2 => std_logic_vector(to_unsigned( 219, 8)),
3 => std_logic_vector(to_unsigned( 194, 8)),
4 => std_logic_vector(to_unsigned( 37, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 198, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 229, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 243, 8)),
12 => std_logic_vector(to_unsigned( 165, 8)),
13 => std_logic_vector(to_unsigned( 228, 8)),
14 => std_logic_vector(to_unsigned( 202, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 403 then count <= 404; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 16, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 74, 8)),
4 => std_logic_vector(to_unsigned( 41, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 52, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 186, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 404 then count <= 405; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 177, 8)),
3 => std_logic_vector(to_unsigned( 19, 8)),
4 => std_logic_vector(to_unsigned( 199, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 215, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 232, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 209, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 405 then count <= 406; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 168, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 157, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 134, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 101, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 203, 8)),
15 => std_logic_vector(to_unsigned( 206, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 406 then count <= 407; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 4, 8)),
5 => std_logic_vector(to_unsigned( 20, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 21, 8)),
10 => std_logic_vector(to_unsigned( 216, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 24, 8)),
13 => std_logic_vector(to_unsigned( 74, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 52, 8)),
16 => std_logic_vector(to_unsigned( 60, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 407 then count <= 408; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 234, 8)),
2 => std_logic_vector(to_unsigned( 207, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 216, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 229, 8)),
7 => std_logic_vector(to_unsigned( 176, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 236, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 1, 8)),
13 => std_logic_vector(to_unsigned( 219, 8)),
14 => std_logic_vector(to_unsigned( 226, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 126, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 209, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 408 then count <= 409; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 32, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 124, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 85, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 21, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 238, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 132, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 409 then count <= 410; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 117, 8)),
5 => std_logic_vector(to_unsigned( 40, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 67, 8)),
15 => std_logic_vector(to_unsigned( 88, 8)),
16 => std_logic_vector(to_unsigned( 83, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 410 then count <= 411; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 235, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 55, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 1, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 186, 8)),
9 => std_logic_vector(to_unsigned( 81, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 33, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 24, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 411 then count <= 412; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 51, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 228, 8)),
11 => std_logic_vector(to_unsigned( 26, 8)),
12 => std_logic_vector(to_unsigned( 218, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 178, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 412 then count <= 413; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 91, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 105, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 249, 8)),
7 => std_logic_vector(to_unsigned( 38, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 60, 8)),
10 => std_logic_vector(to_unsigned( 108, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 33, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 55, 8)),
16 => std_logic_vector(to_unsigned( 213, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 413 then count <= 414; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 87, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 30, 8)),
9 => std_logic_vector(to_unsigned( 126, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 23, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001101
elsif count = 414 then count <= 415; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 19, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 72, 8)),
6 => std_logic_vector(to_unsigned( 216, 8)),
7 => std_logic_vector(to_unsigned( 176, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 59, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 26, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 415 then count <= 416; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 57, 8)),
3 => std_logic_vector(to_unsigned( 232, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 112, 8)),
6 => std_logic_vector(to_unsigned( 71, 8)),
7 => std_logic_vector(to_unsigned( 23, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 141, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 20, 8)),
16 => std_logic_vector(to_unsigned( 253, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 416 then count <= 417; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 18, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 185, 8)),
5 => std_logic_vector(to_unsigned( 12, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 238, 8)),
9 => std_logic_vector(to_unsigned( 78, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 70, 8)),
12 => std_logic_vector(to_unsigned( 177, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 134, 8)),
16 => std_logic_vector(to_unsigned( 105, 8)),
17 => std_logic_vector(to_unsigned( 53, 8)),
18 => std_logic_vector(to_unsigned( 200, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 417 then count <= 418; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 32, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 26, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 107, 8)),
11 => std_logic_vector(to_unsigned( 229, 8)),
12 => std_logic_vector(to_unsigned( 85, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 206, 8)),
16 => std_logic_vector(to_unsigned( 132, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 418 then count <= 419; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 10, 8)),
2 => std_logic_vector(to_unsigned( 3, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 182, 8)),
7 => std_logic_vector(to_unsigned( 240, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 63, 8)),
10 => std_logic_vector(to_unsigned( 165, 8)),
11 => std_logic_vector(to_unsigned( 38, 8)),
12 => std_logic_vector(to_unsigned( 232, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 231, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 419 then count <= 420; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 222, 8)),
4 => std_logic_vector(to_unsigned( 88, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 164, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 208, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 236, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 226, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 420 then count <= 421; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 211, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 50, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 130, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 91, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 421 then count <= 422; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 199, 8)),
2 => std_logic_vector(to_unsigned( 206, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 105, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 85, 8)),
10 => std_logic_vector(to_unsigned( 183, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 237, 8)),
14 => std_logic_vector(to_unsigned( 186, 8)),
15 => std_logic_vector(to_unsigned( 57, 8)),
16 => std_logic_vector(to_unsigned( 245, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110110
elsif count = 422 then count <= 423; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 168, 8)),
2 => std_logic_vector(to_unsigned( 143, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 87, 8)),
11 => std_logic_vector(to_unsigned( 244, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 423 then count <= 424; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 204, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 226, 8)),
5 => std_logic_vector(to_unsigned( 250, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 80, 8)),
10 => std_logic_vector(to_unsigned( 96, 8)),
11 => std_logic_vector(to_unsigned( 173, 8)),
12 => std_logic_vector(to_unsigned( 252, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 216, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 424 then count <= 425; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 243, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 44, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 11, 8)),
8 => std_logic_vector(to_unsigned( 232, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 0, 8)),
16 => std_logic_vector(to_unsigned( 43, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 425 then count <= 426; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 112, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 249, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 246, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 189, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 426 then count <= 427; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 185, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 102, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 63, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 145, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 427 then count <= 428; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 236, 8)),
3 => std_logic_vector(to_unsigned( 231, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 207, 8)),
6 => std_logic_vector(to_unsigned( 34, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 149, 8)),
9 => std_logic_vector(to_unsigned( 0, 8)),
10 => std_logic_vector(to_unsigned( 1, 8)),
11 => std_logic_vector(to_unsigned( 49, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 238, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 79, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 428 then count <= 429; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 111, 8)),
2 => std_logic_vector(to_unsigned( 196, 8)),
3 => std_logic_vector(to_unsigned( 190, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 133, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 198, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 429 then count <= 430; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 12, 8)),
4 => std_logic_vector(to_unsigned( 56, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 135, 8)),
9 => std_logic_vector(to_unsigned( 47, 8)),
10 => std_logic_vector(to_unsigned( 232, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 173, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 177, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 430 then count <= 431; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 139, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 49, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 247, 8)),
7 => std_logic_vector(to_unsigned( 42, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 57, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 218, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010011
elsif count = 431 then count <= 432; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 195, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 231, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 4, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 226, 8)),
14 => std_logic_vector(to_unsigned( 57, 8)),
15 => std_logic_vector(to_unsigned( 68, 8)),
16 => std_logic_vector(to_unsigned( 226, 8)),
17 => std_logic_vector(to_unsigned( 188, 8)),
18 => std_logic_vector(to_unsigned( 52, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 432 then count <= 433; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 25, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 30, 8)),
11 => std_logic_vector(to_unsigned( 3, 8)),
12 => std_logic_vector(to_unsigned( 244, 8)),
13 => std_logic_vector(to_unsigned( 199, 8)),
14 => std_logic_vector(to_unsigned( 186, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 433 then count <= 434; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 204, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 125, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 434 then count <= 435; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 237, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 153, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 247, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 15, 8)),
10 => std_logic_vector(to_unsigned( 252, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 239, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 435 then count <= 436; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 234, 8)),
2 => std_logic_vector(to_unsigned( 206, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 27, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 108, 8)),
8 => std_logic_vector(to_unsigned( 17, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 234, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 44, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 436 then count <= 437; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 247, 8)),
2 => std_logic_vector(to_unsigned( 17, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 215, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 44, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 146, 8)),
15 => std_logic_vector(to_unsigned( 25, 8)),
16 => std_logic_vector(to_unsigned( 59, 8)),
17 => std_logic_vector(to_unsigned( 34, 8)),
18 => std_logic_vector(to_unsigned( 36, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 437 then count <= 438; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 216, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 17, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 138, 8)),
14 => std_logic_vector(to_unsigned( 13, 8)),
15 => std_logic_vector(to_unsigned( 218, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 438 then count <= 439; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 245, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 3, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 245, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 87, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 21, 8)),
14 => std_logic_vector(to_unsigned( 188, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 40, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 439 then count <= 440; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 177, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 230, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 71, 8)),
8 => std_logic_vector(to_unsigned( 186, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 21, 8)),
12 => std_logic_vector(to_unsigned( 84, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 68, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001010
elsif count = 440 then count <= 441; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 205, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 222, 8)),
4 => std_logic_vector(to_unsigned( 75, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 28, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 441 then count <= 442; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 156, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 54, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 229, 8)),
13 => std_logic_vector(to_unsigned( 251, 8)),
14 => std_logic_vector(to_unsigned( 35, 8)),
15 => std_logic_vector(to_unsigned( 74, 8)),
16 => std_logic_vector(to_unsigned( 136, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010101
elsif count = 442 then count <= 443; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 16, 8)),
4 => std_logic_vector(to_unsigned( 228, 8)),
5 => std_logic_vector(to_unsigned( 198, 8)),
6 => std_logic_vector(to_unsigned( 152, 8)),
7 => std_logic_vector(to_unsigned( 213, 8)),
8 => std_logic_vector(to_unsigned( 137, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 199, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 73, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 443 then count <= 444; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 233, 8)),
3 => std_logic_vector(to_unsigned( 13, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 220, 8)),
6 => std_logic_vector(to_unsigned( 26, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 185, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 239, 8)),
11 => std_logic_vector(to_unsigned( 188, 8)),
12 => std_logic_vector(to_unsigned( 193, 8)),
13 => std_logic_vector(to_unsigned( 3, 8)),
14 => std_logic_vector(to_unsigned( 232, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 444 then count <= 445; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 205, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 17, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 35, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 445 then count <= 446; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 242, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 230, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 212, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 231, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 28, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 446 then count <= 447; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 36, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 50, 8)),
6 => std_logic_vector(to_unsigned( 185, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 88, 8)),
13 => std_logic_vector(to_unsigned( 55, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 41, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 447 then count <= 448; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 205, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 20, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 46, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 15, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 221, 8)),
17 => std_logic_vector(to_unsigned( 78, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 448 then count <= 449; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 91, 8)),
2 => std_logic_vector(to_unsigned( 16, 8)),
3 => std_logic_vector(to_unsigned( 204, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 86, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 83, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 237, 8)),
14 => std_logic_vector(to_unsigned( 185, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 449 then count <= 450; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 197, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 156, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 163, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 450 then count <= 451; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 226, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 241, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 217, 8)),
8 => std_logic_vector(to_unsigned( 57, 8)),
9 => std_logic_vector(to_unsigned( 199, 8)),
10 => std_logic_vector(to_unsigned( 59, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 121, 8)),
17 => std_logic_vector(to_unsigned( 209, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 451 then count <= 452; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 141, 8)),
3 => std_logic_vector(to_unsigned( 45, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 231, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 236, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 452 then count <= 453; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 104, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 253, 8)),
8 => std_logic_vector(to_unsigned( 54, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 129, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 453 then count <= 454; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 21, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 243, 8)),
5 => std_logic_vector(to_unsigned( 61, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 253, 8)),
11 => std_logic_vector(to_unsigned( 249, 8)),
12 => std_logic_vector(to_unsigned( 233, 8)),
13 => std_logic_vector(to_unsigned( 55, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 46, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 48, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 454 then count <= 455; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 78, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 55, 8)),
4 => std_logic_vector(to_unsigned( 8, 8)),
5 => std_logic_vector(to_unsigned( 119, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 57, 8)),
9 => std_logic_vector(to_unsigned( 33, 8)),
10 => std_logic_vector(to_unsigned( 28, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 38, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 246, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 168, 8)),
17 => std_logic_vector(to_unsigned( 54, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 455 then count <= 456; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 89, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 207, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 78, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 49, 8)),
16 => std_logic_vector(to_unsigned( 64, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 456 then count <= 457; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 173, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 238, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 96, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 37, 8)),
16 => std_logic_vector(to_unsigned( 214, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 457 then count <= 458; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 67, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 28, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 127, 8)),
9 => std_logic_vector(to_unsigned( 45, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 16, 8)),
12 => std_logic_vector(to_unsigned( 90, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 50, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 458 then count <= 459; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 214, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 66, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 92, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 123, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 459 then count <= 460; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 254, 8)),
2 => std_logic_vector(to_unsigned( 198, 8)),
3 => std_logic_vector(to_unsigned( 109, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 88, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 217, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 200, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101100
elsif count = 460 then count <= 461; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 7, 8)),
6 => std_logic_vector(to_unsigned( 20, 8)),
7 => std_logic_vector(to_unsigned( 7, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 96, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110010
elsif count = 461 then count <= 462; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 105, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 236, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 91, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 212, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 165, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 462 then count <= 463; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 33, 8)),
2 => std_logic_vector(to_unsigned( 202, 8)),
3 => std_logic_vector(to_unsigned( 199, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 214, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 246, 8)),
12 => std_logic_vector(to_unsigned( 77, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 226, 8)),
17 => std_logic_vector(to_unsigned( 215, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 463 then count <= 464; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 47, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010110
elsif count = 464 then count <= 465; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 21, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 189, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 161, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 135, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 78, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 465 then count <= 466; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 100, 8)),
4 => std_logic_vector(to_unsigned( 112, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 27, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 134, 8)),
16 => std_logic_vector(to_unsigned( 26, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 466 then count <= 467; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 84, 8)),
4 => std_logic_vector(to_unsigned( 215, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 220, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 4, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 467 then count <= 468; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 43, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 77, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 101, 8)),
8 => std_logic_vector(to_unsigned( 109, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 54, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 36, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 468 then count <= 469; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 33, 8)),
6 => std_logic_vector(to_unsigned( 89, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 60, 8)),
9 => std_logic_vector(to_unsigned( 184, 8)),
10 => std_logic_vector(to_unsigned( 173, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 43, 8)),
14 => std_logic_vector(to_unsigned( 181, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 469 then count <= 470; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 3, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 218, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 231, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 242, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 147, 8)),
12 => std_logic_vector(to_unsigned( 168, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 214, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 239, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 185, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 470 then count <= 471; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 226, 8)),
5 => std_logic_vector(to_unsigned( 197, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 154, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 95, 8)),
14 => std_logic_vector(to_unsigned( 203, 8)),
15 => std_logic_vector(to_unsigned( 172, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 471 then count <= 472; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 193, 8)),
7 => std_logic_vector(to_unsigned( 11, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 119, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 196, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 113, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110110
elsif count = 472 then count <= 473; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 251, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 80, 8)),
4 => std_logic_vector(to_unsigned( 30, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 207, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 20, 8)),
12 => std_logic_vector(to_unsigned( 177, 8)),
13 => std_logic_vector(to_unsigned( 31, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 33, 8)),
16 => std_logic_vector(to_unsigned( 0, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 473 then count <= 474; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 32, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 239, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 49, 8)),
12 => std_logic_vector(to_unsigned( 41, 8)),
13 => std_logic_vector(to_unsigned( 35, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 52, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 474 then count <= 475; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 12, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 88, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 132, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 145, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 54, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 90, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 475 then count <= 476; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 130, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 3, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 190, 8)),
6 => std_logic_vector(to_unsigned( 236, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 60, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 476 then count <= 477; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 249, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 39, 8)),
7 => std_logic_vector(to_unsigned( 27, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 63, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 209, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110011
elsif count = 477 then count <= 478; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 232, 8)),
12 => std_logic_vector(to_unsigned( 154, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 147, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 478 then count <= 479; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 32, 8)),
2 => std_logic_vector(to_unsigned( 37, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 227, 8)),
6 => std_logic_vector(to_unsigned( 207, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 162, 8)),
11 => std_logic_vector(to_unsigned( 34, 8)),
12 => std_logic_vector(to_unsigned( 41, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 22, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 38, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 479 then count <= 480; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 75, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 169, 8)),
9 => std_logic_vector(to_unsigned( 212, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 168, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 188, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 480 then count <= 481; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 20, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 248, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 170, 8)),
6 => std_logic_vector(to_unsigned( 94, 8)),
7 => std_logic_vector(to_unsigned( 147, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 147, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 481 then count <= 482; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 198, 8)),
3 => std_logic_vector(to_unsigned( 149, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 59, 8)),
9 => std_logic_vector(to_unsigned( 98, 8)),
10 => std_logic_vector(to_unsigned( 166, 8)),
11 => std_logic_vector(to_unsigned( 55, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 51, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110101
elsif count = 482 then count <= 483; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 22, 8)),
3 => std_logic_vector(to_unsigned( 30, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 40, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 230, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 47, 8)),
14 => std_logic_vector(to_unsigned( 52, 8)),
15 => std_logic_vector(to_unsigned( 81, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 91, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 483 then count <= 484; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 16, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 46, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 247, 8)),
8 => std_logic_vector(to_unsigned( 182, 8)),
9 => std_logic_vector(to_unsigned( 107, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 243, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 51, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 484 then count <= 485; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 222, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 116, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 15, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 219, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 251, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 192, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 212, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 485 then count <= 486; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 116, 8)),
2 => std_logic_vector(to_unsigned( 193, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 251, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 192, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 116, 8)),
15 => std_logic_vector(to_unsigned( 177, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 76, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 486 then count <= 487; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 22, 8)),
2 => std_logic_vector(to_unsigned( 196, 8)),
3 => std_logic_vector(to_unsigned( 23, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 19, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 197, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 68, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 487 then count <= 488; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 243, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 26, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 218, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 179, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 250, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 205, 8)),
18 => std_logic_vector(to_unsigned( 181, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 488 then count <= 489; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 9, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 165, 8)),
4 => std_logic_vector(to_unsigned( 32, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 6, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 56, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 165, 8)),
15 => std_logic_vector(to_unsigned( 143, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 489 then count <= 490; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 12, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 184, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 5, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 69, 8)),
14 => std_logic_vector(to_unsigned( 44, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 145, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 40, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 490 then count <= 491; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 42, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 33, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 163, 8)),
14 => std_logic_vector(to_unsigned( 6, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 491 then count <= 492; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 229, 8)),
7 => std_logic_vector(to_unsigned( 0, 8)),
8 => std_logic_vector(to_unsigned( 8, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 28, 8)),
12 => std_logic_vector(to_unsigned( 63, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 198, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 229, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 198, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 492 then count <= 493; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 88, 8)),
3 => std_logic_vector(to_unsigned( 34, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 49, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 4, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 35, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 493 then count <= 494; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 171, 8)),
2 => std_logic_vector(to_unsigned( 130, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 77, 8)),
5 => std_logic_vector(to_unsigned( 77, 8)),
6 => std_logic_vector(to_unsigned( 29, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 192, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 87, 8)),
14 => std_logic_vector(to_unsigned( 19, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 53, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 494 then count <= 495; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 4, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 68, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 179, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 495 then count <= 496; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 71, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 30, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 21, 8)),
6 => std_logic_vector(to_unsigned( 235, 8)),
7 => std_logic_vector(to_unsigned( 84, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 14, 8)),
12 => std_logic_vector(to_unsigned( 145, 8)),
13 => std_logic_vector(to_unsigned( 22, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 194, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 55, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 496 then count <= 497; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 152, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 200, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 230, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 240, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 232, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 172, 8)),
16 => std_logic_vector(to_unsigned( 60, 8)),
17 => std_logic_vector(to_unsigned( 196, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 497 then count <= 498; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 81, 8)),
2 => std_logic_vector(to_unsigned( 156, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 116, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 41, 8)),
9 => std_logic_vector(to_unsigned( 222, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 88, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 498 then count <= 499; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 30, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 139, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 24, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 221, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 499 then count <= 500; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 226, 8)),
2 => std_logic_vector(to_unsigned( 82, 8)),
3 => std_logic_vector(to_unsigned( 209, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 184, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 212, 8)),
10 => std_logic_vector(to_unsigned( 68, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 84, 8)),
13 => std_logic_vector(to_unsigned( 212, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 233, 8)),
16 => std_logic_vector(to_unsigned( 89, 8)),
17 => std_logic_vector(to_unsigned( 203, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 500 then count <= 501; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 171, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 181, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 200, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 187, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 501 then count <= 502; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 35, 8)),
2 => std_logic_vector(to_unsigned( 121, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 204, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 39, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 502 then count <= 503; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 177, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 15, 8)),
15 => std_logic_vector(to_unsigned( 127, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100110
elsif count = 503 then count <= 504; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 158, 8)),
3 => std_logic_vector(to_unsigned( 240, 8)),
4 => std_logic_vector(to_unsigned( 208, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 135, 8)),
9 => std_logic_vector(to_unsigned( 182, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 207, 8)),
12 => std_logic_vector(to_unsigned( 145, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 147, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 504 then count <= 505; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 141, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 38, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 101, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 47, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 87, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 505 then count <= 506; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 142, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 225, 8)),
8 => std_logic_vector(to_unsigned( 149, 8)),
9 => std_logic_vector(to_unsigned( 16, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 179, 8)),
14 => std_logic_vector(to_unsigned( 195, 8)),
15 => std_logic_vector(to_unsigned( 74, 8)),
16 => std_logic_vector(to_unsigned( 234, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 506 then count <= 507; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 159, 8)),
6 => std_logic_vector(to_unsigned( 35, 8)),
7 => std_logic_vector(to_unsigned( 23, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 60, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 1, 8)),
16 => std_logic_vector(to_unsigned( 245, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 507 then count <= 508; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 254, 8)),
4 => std_logic_vector(to_unsigned( 184, 8)),
5 => std_logic_vector(to_unsigned( 100, 8)),
6 => std_logic_vector(to_unsigned( 87, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 140, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 90, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 508 then count <= 509; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 81, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 99, 8)),
5 => std_logic_vector(to_unsigned( 55, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 208, 8)),
8 => std_logic_vector(to_unsigned( 6, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 16, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 86, 8)),
13 => std_logic_vector(to_unsigned( 48, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 63, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 509 then count <= 510; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 204, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 255, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 63, 8)),
9 => std_logic_vector(to_unsigned( 198, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 236, 8)),
14 => std_logic_vector(to_unsigned( 180, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011001
elsif count = 510 then count <= 511; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 209, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 178, 8)),
5 => std_logic_vector(to_unsigned( 220, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 181, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 150, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 241, 8)),
14 => std_logic_vector(to_unsigned( 244, 8)),
15 => std_logic_vector(to_unsigned( 2, 8)),
16 => std_logic_vector(to_unsigned( 246, 8)),
17 => std_logic_vector(to_unsigned( 189, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 511 then count <= 512; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 249, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 147, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 58, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 512 then count <= 513; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 112, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 242, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 21, 8)),
13 => std_logic_vector(to_unsigned( 224, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 177, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 513 then count <= 514; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 17, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 91, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 514 then count <= 515; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 81, 8)),
2 => std_logic_vector(to_unsigned( 31, 8)),
3 => std_logic_vector(to_unsigned( 113, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 224, 8)),
7 => std_logic_vector(to_unsigned( 60, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 29, 8)),
11 => std_logic_vector(to_unsigned( 36, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 133, 8)),
14 => std_logic_vector(to_unsigned( 79, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 515 then count <= 516; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 201, 8)),
3 => std_logic_vector(to_unsigned( 68, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 103, 8)),
8 => std_logic_vector(to_unsigned( 197, 8)),
9 => std_logic_vector(to_unsigned( 57, 8)),
10 => std_logic_vector(to_unsigned( 2, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 218, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 6, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 516 then count <= 517; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 180, 8)),
2 => std_logic_vector(to_unsigned( 76, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 72, 8)),
12 => std_logic_vector(to_unsigned( 227, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 62, 8)),
15 => std_logic_vector(to_unsigned( 164, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 517 then count <= 518; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 242, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 237, 8)),
4 => std_logic_vector(to_unsigned( 116, 8)),
5 => std_logic_vector(to_unsigned( 9, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 100, 8)),
9 => std_logic_vector(to_unsigned( 45, 8)),
10 => std_logic_vector(to_unsigned( 163, 8)),
11 => std_logic_vector(to_unsigned( 60, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 188, 8)),
15 => std_logic_vector(to_unsigned( 38, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 518 then count <= 519; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 160, 8)),
3 => std_logic_vector(to_unsigned( 74, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 2, 8)),
6 => std_logic_vector(to_unsigned( 182, 8)),
7 => std_logic_vector(to_unsigned( 147, 8)),
8 => std_logic_vector(to_unsigned( 241, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 99, 8)),
16 => std_logic_vector(to_unsigned( 221, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 519 then count <= 520; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 68, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 224, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 220, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 241, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 43, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 197, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 520 then count <= 521; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 204, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 212, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 116, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 11, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110010
elsif count = 521 then count <= 522; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 177, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 110, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 191, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 11, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 522 then count <= 523; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 227, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 233, 8)),
4 => std_logic_vector(to_unsigned( 108, 8)),
5 => std_logic_vector(to_unsigned( 192, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 65, 8)),
12 => std_logic_vector(to_unsigned( 187, 8)),
13 => std_logic_vector(to_unsigned( 240, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 229, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 202, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 523 then count <= 524; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 44, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 38, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 9, 8)),
9 => std_logic_vector(to_unsigned( 243, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 55, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 79, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 19, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 524 then count <= 525; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 79, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 109, 8)),
6 => std_logic_vector(to_unsigned( 233, 8)),
7 => std_logic_vector(to_unsigned( 219, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 228, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 223, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 54, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 525 then count <= 526; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 215, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 204, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 16, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 55, 8)),
11 => std_logic_vector(to_unsigned( 12, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 229, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 526 then count <= 527; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 221, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 215, 8)),
8 => std_logic_vector(to_unsigned( 93, 8)),
9 => std_logic_vector(to_unsigned( 138, 8)),
10 => std_logic_vector(to_unsigned( 182, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 100, 8)),
15 => std_logic_vector(to_unsigned( 234, 8)),
16 => std_logic_vector(to_unsigned( 1, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00001111
elsif count = 527 then count <= 528; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 61, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 49, 8)),
5 => std_logic_vector(to_unsigned( 39, 8)),
6 => std_logic_vector(to_unsigned( 173, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 150, 8)),
12 => std_logic_vector(to_unsigned( 193, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 73, 8)),
17 => std_logic_vector(to_unsigned( 64, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 528 then count <= 529; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 35, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 238, 8)),
7 => std_logic_vector(to_unsigned( 212, 8)),
8 => std_logic_vector(to_unsigned( 245, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 175, 8)),
14 => std_logic_vector(to_unsigned( 231, 8)),
15 => std_logic_vector(to_unsigned( 238, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 529 then count <= 530; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 232, 8)),
2 => std_logic_vector(to_unsigned( 241, 8)),
3 => std_logic_vector(to_unsigned( 239, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 195, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 191, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 132, 8)),
12 => std_logic_vector(to_unsigned( 191, 8)),
13 => std_logic_vector(to_unsigned( 249, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 530 then count <= 531; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 200, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 165, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 240, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 5, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 230, 8)),
12 => std_logic_vector(to_unsigned( 44, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 223, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 531 then count <= 532; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 86, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 22, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 532 then count <= 533; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 247, 8)),
4 => std_logic_vector(to_unsigned( 99, 8)),
5 => std_logic_vector(to_unsigned( 159, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 86, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 32, 8)),
14 => std_logic_vector(to_unsigned( 188, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 533 then count <= 534; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 76, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 237, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 54, 8)),
9 => std_logic_vector(to_unsigned( 222, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 156, 8)),
12 => std_logic_vector(to_unsigned( 68, 8)),
13 => std_logic_vector(to_unsigned( 53, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 534 then count <= 535; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 225, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 174, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 213, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 84, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 224, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 221, 8)),
15 => std_logic_vector(to_unsigned( 209, 8)),
16 => std_logic_vector(to_unsigned( 205, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 535 then count <= 536; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 195, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 229, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 205, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 63, 8)),
9 => std_logic_vector(to_unsigned( 202, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 189, 8)),
13 => std_logic_vector(to_unsigned( 64, 8)),
14 => std_logic_vector(to_unsigned( 140, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 32, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 61, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 536 then count <= 537; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 16, 8)),
2 => std_logic_vector(to_unsigned( 2, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 249, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 44, 8)),
8 => std_logic_vector(to_unsigned( 212, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 40, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 183, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 537 then count <= 538; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 199, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 232, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 237, 8)),
8 => std_logic_vector(to_unsigned( 97, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 71, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 51, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 245, 8)),
16 => std_logic_vector(to_unsigned( 89, 8)),
17 => std_logic_vector(to_unsigned( 217, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 538 then count <= 539; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 197, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 252, 8)),
7 => std_logic_vector(to_unsigned( 210, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 115, 8)),
11 => std_logic_vector(to_unsigned( 153, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 63, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 539 then count <= 540; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 232, 8)),
7 => std_logic_vector(to_unsigned( 221, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 146, 8)),
10 => std_logic_vector(to_unsigned( 184, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 175, 8)),
14 => std_logic_vector(to_unsigned( 213, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 247, 8)),
17 => std_logic_vector(to_unsigned( 190, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 540 then count <= 541; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 111, 8)),
2 => std_logic_vector(to_unsigned( 5, 8)),
3 => std_logic_vector(to_unsigned( 213, 8)),
4 => std_logic_vector(to_unsigned( 88, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 26, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 142, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 16, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101010
elsif count = 541 then count <= 542; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 222, 8)),
4 => std_logic_vector(to_unsigned( 8, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 24, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 227, 8)),
12 => std_logic_vector(to_unsigned( 160, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 542 then count <= 543; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 35, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 90, 8)),
4 => std_logic_vector(to_unsigned( 20, 8)),
5 => std_logic_vector(to_unsigned( 173, 8)),
6 => std_logic_vector(to_unsigned( 14, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 63, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 39, 8)),
11 => std_logic_vector(to_unsigned( 66, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 147, 8)),
15 => std_logic_vector(to_unsigned( 232, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 52, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111010
elsif count = 543 then count <= 544; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 20, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 136, 8)),
10 => std_logic_vector(to_unsigned( 95, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 150, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 74, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 62, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 544 then count <= 545; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 62, 8)),
2 => std_logic_vector(to_unsigned( 235, 8)),
3 => std_logic_vector(to_unsigned( 222, 8)),
4 => std_logic_vector(to_unsigned( 235, 8)),
5 => std_logic_vector(to_unsigned( 219, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 239, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 21, 8)),
14 => std_logic_vector(to_unsigned( 226, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 545 then count <= 546; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 229, 8)),
2 => std_logic_vector(to_unsigned( 194, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 230, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 104, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 236, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 157, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 546 then count <= 547; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 45, 8)),
4 => std_logic_vector(to_unsigned( 207, 8)),
5 => std_logic_vector(to_unsigned( 115, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 63, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 12, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 547 then count <= 548; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 43, 8)),
2 => std_logic_vector(to_unsigned( 236, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 51, 8)),
6 => std_logic_vector(to_unsigned( 94, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 97, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 188, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 44, 8)),
15 => std_logic_vector(to_unsigned( 223, 8)),
16 => std_logic_vector(to_unsigned( 235, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 548 then count <= 549; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 208, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 17, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 155, 8)),
9 => std_logic_vector(to_unsigned( 181, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 229, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 182, 8)),
16 => std_logic_vector(to_unsigned( 233, 8)),
17 => std_logic_vector(to_unsigned( 202, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 549 then count <= 550; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 204, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 213, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 240, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 10, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 79, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 192, 8)),
13 => std_logic_vector(to_unsigned( 94, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 550 then count <= 551; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 143, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 89, 8)),
5 => std_logic_vector(to_unsigned( 181, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 110, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 249, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 222, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010011
elsif count = 551 then count <= 552; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 74, 8)),
4 => std_logic_vector(to_unsigned( 61, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 85, 8)),
13 => std_logic_vector(to_unsigned( 247, 8)),
14 => std_logic_vector(to_unsigned( 234, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 50, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 552 then count <= 553; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 81, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 151, 8)),
4 => std_logic_vector(to_unsigned( 55, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 123, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 28, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 35, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 244, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 553 then count <= 554; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 148, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 17, 8)),
11 => std_logic_vector(to_unsigned( 232, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 59, 8)),
14 => std_logic_vector(to_unsigned( 226, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 554 then count <= 555; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 84, 8)),
3 => std_logic_vector(to_unsigned( 50, 8)),
4 => std_logic_vector(to_unsigned( 18, 8)),
5 => std_logic_vector(to_unsigned( 51, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 16, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 63, 8)),
11 => std_logic_vector(to_unsigned( 18, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 53, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 48, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 555 then count <= 556; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 241, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 21, 8)),
5 => std_logic_vector(to_unsigned( 254, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 72, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 38, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 7, 8)),
15 => std_logic_vector(to_unsigned( 128, 8)),
16 => std_logic_vector(to_unsigned( 185, 8)),
17 => std_logic_vector(to_unsigned( 206, 8)),
18 => std_logic_vector(to_unsigned( 51, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00100111
elsif count = 556 then count <= 557; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 234, 8)),
2 => std_logic_vector(to_unsigned( 145, 8)),
3 => std_logic_vector(to_unsigned( 41, 8)),
4 => std_logic_vector(to_unsigned( 219, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 221, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 40, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 223, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 207, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 557 then count <= 558; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 37, 8)),
4 => std_logic_vector(to_unsigned( 224, 8)),
5 => std_logic_vector(to_unsigned( 149, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 184, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 203, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 558 then count <= 559; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 129, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 4, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 139, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 95, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 47, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 128, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 559 then count <= 560; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 128, 8)),
2 => std_logic_vector(to_unsigned( 0, 8)),
3 => std_logic_vector(to_unsigned( 84, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 58, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 560 then count <= 561; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 205, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 142, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 244, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 139, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010110
elsif count = 561 then count <= 562; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 165, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 140, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 218, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 222, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 68, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 562 then count <= 563; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 221, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 170, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 160, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 24, 8)),
9 => std_logic_vector(to_unsigned( 233, 8)),
10 => std_logic_vector(to_unsigned( 36, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 253, 8)),
16 => std_logic_vector(to_unsigned( 51, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00100111
elsif count = 563 then count <= 564; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 112, 8)),
3 => std_logic_vector(to_unsigned( 80, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 99, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 236, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 564 then count <= 565; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 9, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 95, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 213, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 565 then count <= 566; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 121, 8)),
3 => std_logic_vector(to_unsigned( 208, 8)),
4 => std_logic_vector(to_unsigned( 117, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 241, 8)),
8 => std_logic_vector(to_unsigned( 169, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 150, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 566 then count <= 567; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 230, 8)),
4 => std_logic_vector(to_unsigned( 200, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 215, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 10, 8)),
14 => std_logic_vector(to_unsigned( 128, 8)),
15 => std_logic_vector(to_unsigned( 147, 8)),
16 => std_logic_vector(to_unsigned( 225, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 200, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 567 then count <= 568; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 0, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 98, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 238, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 51, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 568 then count <= 569; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 40, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 132, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 105, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 569 then count <= 570; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 155, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 181, 8)),
5 => std_logic_vector(to_unsigned( 164, 8)),
6 => std_logic_vector(to_unsigned( 137, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 231, 8)),
13 => std_logic_vector(to_unsigned( 202, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 92, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 570 then count <= 571; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 32, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 239, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 217, 8)),
8 => std_logic_vector(to_unsigned( 16, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 122, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 141, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100100
elsif count = 571 then count <= 572; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 24, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 229, 8)),
6 => std_logic_vector(to_unsigned( 12, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 251, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 236, 8)),
13 => std_logic_vector(to_unsigned( 45, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 206, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111010
elsif count = 572 then count <= 573; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 192, 8)),
12 => std_logic_vector(to_unsigned( 1, 8)),
13 => std_logic_vector(to_unsigned( 208, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 573 then count <= 574; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 31, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 156, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 203, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 18, 8)),
12 => std_logic_vector(to_unsigned( 238, 8)),
13 => std_logic_vector(to_unsigned( 201, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 211, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 184, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 574 then count <= 575; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 226, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 30, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 3, 8)),
11 => std_logic_vector(to_unsigned( 66, 8)),
12 => std_logic_vector(to_unsigned( 1, 8)),
13 => std_logic_vector(to_unsigned( 100, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 21, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 575 then count <= 576; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 185, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 35, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 67, 8)),
7 => std_logic_vector(to_unsigned( 244, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 210, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 34, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 195, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 576 then count <= 577; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 22, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 101, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 220, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 577 then count <= 578; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 62, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 249, 8)),
6 => std_logic_vector(to_unsigned( 74, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 76, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 254, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 123, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001011
elsif count = 578 then count <= 579; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 181, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 243, 8)),
6 => std_logic_vector(to_unsigned( 235, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 29, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 1, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 211, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 208, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 579 then count <= 580; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 198, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 77, 8)),
9 => std_logic_vector(to_unsigned( 118, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 32, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 580 then count <= 581; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 28, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 2, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 54, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 46, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 581 then count <= 582; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 3, 8)),
5 => std_logic_vector(to_unsigned( 220, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 170, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 250, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 216, 8)),
14 => std_logic_vector(to_unsigned( 185, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 131, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 582 then count <= 583; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 16, 8)),
5 => std_logic_vector(to_unsigned( 207, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 32, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 18, 8)),
15 => std_logic_vector(to_unsigned( 71, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 29, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 583 then count <= 584; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 70, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 210, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 254, 8)),
9 => std_logic_vector(to_unsigned( 218, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 35, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 59, 8)),
15 => std_logic_vector(to_unsigned( 209, 8)),
16 => std_logic_vector(to_unsigned( 245, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 584 then count <= 585; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 54, 8)),
3 => std_logic_vector(to_unsigned( 154, 8)),
4 => std_logic_vector(to_unsigned( 49, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 66, 8)),
9 => std_logic_vector(to_unsigned( 78, 8)),
10 => std_logic_vector(to_unsigned( 95, 8)),
11 => std_logic_vector(to_unsigned( 193, 8)),
12 => std_logic_vector(to_unsigned( 88, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 585 then count <= 586; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 233, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 212, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 136, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 22, 8)),
12 => std_logic_vector(to_unsigned( 24, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 141, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 168, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 586 then count <= 587; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 33, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 155, 8)),
5 => std_logic_vector(to_unsigned( 11, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 239, 8)),
8 => std_logic_vector(to_unsigned( 226, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 36, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 26, 8)),
13 => std_logic_vector(to_unsigned( 100, 8)),
14 => std_logic_vector(to_unsigned( 80, 8)),
15 => std_logic_vector(to_unsigned( 80, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 53, 8)),
18 => std_logic_vector(to_unsigned( 60, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110101
elsif count = 587 then count <= 588; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 30, 8)),
2 => std_logic_vector(to_unsigned( 190, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 166, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 198, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 235, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 48, 8)),
12 => std_logic_vector(to_unsigned( 218, 8)),
13 => std_logic_vector(to_unsigned( 7, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 74, 8)),
16 => std_logic_vector(to_unsigned( 48, 8)),
17 => std_logic_vector(to_unsigned( 73, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 588 then count <= 589; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 60, 8)),
3 => std_logic_vector(to_unsigned( 129, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 2, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 589 then count <= 590; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 155, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 12, 8)),
6 => std_logic_vector(to_unsigned( 245, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 92, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 10, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 133, 8)),
14 => std_logic_vector(to_unsigned( 17, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 15, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 590 then count <= 591; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 11, 8)),
2 => std_logic_vector(to_unsigned( 254, 8)),
3 => std_logic_vector(to_unsigned( 234, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 240, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 139, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011000
elsif count = 591 then count <= 592; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 125, 8)),
3 => std_logic_vector(to_unsigned( 254, 8)),
4 => std_logic_vector(to_unsigned( 228, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 71, 8)),
11 => std_logic_vector(to_unsigned( 62, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 44, 8)),
14 => std_logic_vector(to_unsigned( 216, 8)),
15 => std_logic_vector(to_unsigned( 251, 8)),
16 => std_logic_vector(to_unsigned( 141, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 592 then count <= 593; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 253, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 211, 8)),
8 => std_logic_vector(to_unsigned( 26, 8)),
9 => std_logic_vector(to_unsigned( 176, 8)),
10 => std_logic_vector(to_unsigned( 76, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 593 then count <= 594; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 4, 8)),
2 => std_logic_vector(to_unsigned( 234, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 184, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 186, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 95, 8)),
12 => std_logic_vector(to_unsigned( 53, 8)),
13 => std_logic_vector(to_unsigned( 95, 8)),
14 => std_logic_vector(to_unsigned( 234, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 204, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011010
elsif count = 594 then count <= 595; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 95, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 71, 8)),
5 => std_logic_vector(to_unsigned( 58, 8)),
6 => std_logic_vector(to_unsigned( 11, 8)),
7 => std_logic_vector(to_unsigned( 103, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 119, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 139, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 595 then count <= 596; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 217, 8)),
5 => std_logic_vector(to_unsigned( 189, 8)),
6 => std_logic_vector(to_unsigned( 33, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 66, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 186, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 596 then count <= 597; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 235, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 174, 8)),
4 => std_logic_vector(to_unsigned( 208, 8)),
5 => std_logic_vector(to_unsigned( 221, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 213, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 0, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110110
elsif count = 597 then count <= 598; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 246, 8)),
2 => std_logic_vector(to_unsigned( 158, 8)),
3 => std_logic_vector(to_unsigned( 239, 8)),
4 => std_logic_vector(to_unsigned( 248, 8)),
5 => std_logic_vector(to_unsigned( 225, 8)),
6 => std_logic_vector(to_unsigned( 137, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 212, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 244, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 147, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 598 then count <= 599; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 39, 8)),
6 => std_logic_vector(to_unsigned( 19, 8)),
7 => std_logic_vector(to_unsigned( 132, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 148, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 244, 8)),
12 => std_logic_vector(to_unsigned( 187, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 194, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 599 then count <= 600; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 142, 8)),
3 => std_logic_vector(to_unsigned( 29, 8)),
4 => std_logic_vector(to_unsigned( 158, 8)),
5 => std_logic_vector(to_unsigned( 104, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 23, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 18, 8)),
11 => std_logic_vector(to_unsigned( 48, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 12, 8)),
15 => std_logic_vector(to_unsigned( 47, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 81, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 600 then count <= 601; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 166, 8)),
8 => std_logic_vector(to_unsigned( 55, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 11, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 243, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 202, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 141, 8)),
17 => std_logic_vector(to_unsigned( 181, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 601 then count <= 602; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 179, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 222, 8)),
5 => std_logic_vector(to_unsigned( 90, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 161, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 53, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 249, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 602 then count <= 603; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 91, 8)),
3 => std_logic_vector(to_unsigned( 47, 8)),
4 => std_logic_vector(to_unsigned( 34, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 131, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 212, 8)),
11 => std_logic_vector(to_unsigned( 223, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 224, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 10, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 603 then count <= 604; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 79, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 222, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 232, 8)),
7 => std_logic_vector(to_unsigned( 212, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 246, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 245, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 214, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 604 then count <= 605; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 37, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 47, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 85, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 65, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 13, 8)),
16 => std_logic_vector(to_unsigned( 249, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 605 then count <= 606; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 26, 8)),
3 => std_logic_vector(to_unsigned( 29, 8)),
4 => std_logic_vector(to_unsigned( 217, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 182, 8)),
13 => std_logic_vector(to_unsigned( 79, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 606 then count <= 607; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 180, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 156, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 227, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 141, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 244, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 251, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 607 then count <= 608; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 233, 8)),
2 => std_logic_vector(to_unsigned( 179, 8)),
3 => std_logic_vector(to_unsigned( 246, 8)),
4 => std_logic_vector(to_unsigned( 166, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 199, 8)),
8 => std_logic_vector(to_unsigned( 213, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 216, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 247, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 608 then count <= 609; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 27, 8)),
5 => std_logic_vector(to_unsigned( 100, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 212, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 223, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 609 then count <= 610; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 48, 8)),
6 => std_logic_vector(to_unsigned( 79, 8)),
7 => std_logic_vector(to_unsigned( 189, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 181, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 45, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 78, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 610 then count <= 611; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 216, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 179, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 94, 8)),
8 => std_logic_vector(to_unsigned( 242, 8)),
9 => std_logic_vector(to_unsigned( 89, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 611 then count <= 612; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 186, 8)),
2 => std_logic_vector(to_unsigned( 152, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 91, 8)),
6 => std_logic_vector(to_unsigned( 159, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 64, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 33, 8)),
13 => std_logic_vector(to_unsigned( 94, 8)),
14 => std_logic_vector(to_unsigned( 6, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 131, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 612 then count <= 613; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 226, 8)),
2 => std_logic_vector(to_unsigned( 248, 8)),
3 => std_logic_vector(to_unsigned( 216, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 228, 8)),
9 => std_logic_vector(to_unsigned( 242, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 176, 8)),
12 => std_logic_vector(to_unsigned( 219, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 221, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 613 then count <= 614; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 216, 8)),
2 => std_logic_vector(to_unsigned( 21, 8)),
3 => std_logic_vector(to_unsigned( 169, 8)),
4 => std_logic_vector(to_unsigned( 88, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 104, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 200, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 216, 8)),
16 => std_logic_vector(to_unsigned( 1, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 614 then count <= 615; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 155, 8)),
2 => std_logic_vector(to_unsigned( 28, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 164, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 103, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 189, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 235, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 615 then count <= 616; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 111, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 65, 8)),
4 => std_logic_vector(to_unsigned( 195, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 209, 8)),
7 => std_logic_vector(to_unsigned( 116, 8)),
8 => std_logic_vector(to_unsigned( 214, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 199, 8)),
13 => std_logic_vector(to_unsigned( 208, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 201, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 616 then count <= 617; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 214, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 224, 8)),
11 => std_logic_vector(to_unsigned( 229, 8)),
12 => std_logic_vector(to_unsigned( 151, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 617 then count <= 618; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 85, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 73, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 195, 8)),
7 => std_logic_vector(to_unsigned( 1, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 86, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 205, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 618 then count <= 619; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 166, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 32, 8)),
8 => std_logic_vector(to_unsigned( 63, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 29, 8)),
13 => std_logic_vector(to_unsigned( 176, 8)),
14 => std_logic_vector(to_unsigned( 145, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111010
elsif count = 619 then count <= 620; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 146, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 35, 8)),
4 => std_logic_vector(to_unsigned( 37, 8)),
5 => std_logic_vector(to_unsigned( 40, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 104, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 27, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 95, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 620 then count <= 621; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 141, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 251, 8)),
5 => std_logic_vector(to_unsigned( 173, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 47, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 141, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 246, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 154, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010101
elsif count = 621 then count <= 622; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 128, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 218, 8)),
4 => std_logic_vector(to_unsigned( 247, 8)),
5 => std_logic_vector(to_unsigned( 216, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 181, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 159, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 622 then count <= 623; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 95, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 174, 8)),
4 => std_logic_vector(to_unsigned( 178, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 236, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 208, 8)),
15 => std_logic_vector(to_unsigned( 227, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010011
elsif count = 623 then count <= 624; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 127, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 21, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 217, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 0, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 624 then count <= 625; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 231, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 177, 8)),
5 => std_logic_vector(to_unsigned( 164, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 69, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 19, 8)),
12 => std_logic_vector(to_unsigned( 10, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 625 then count <= 626; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 77, 8)),
5 => std_logic_vector(to_unsigned( 78, 8)),
6 => std_logic_vector(to_unsigned( 184, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 112, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 108, 8)),
11 => std_logic_vector(to_unsigned( 18, 8)),
12 => std_logic_vector(to_unsigned( 186, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 252, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 626 then count <= 627; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 207, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 220, 8)),
8 => std_logic_vector(to_unsigned( 74, 8)),
9 => std_logic_vector(to_unsigned( 11, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 627 then count <= 628; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 182, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 166, 8)),
5 => std_logic_vector(to_unsigned( 1, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 185, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 202, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 628 then count <= 629; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 1, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 34, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 192, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 29, 8)),
16 => std_logic_vector(to_unsigned( 132, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 629 then count <= 630; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 67, 8)),
2 => std_logic_vector(to_unsigned( 227, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 149, 8)),
6 => std_logic_vector(to_unsigned( 70, 8)),
7 => std_logic_vector(to_unsigned( 188, 8)),
8 => std_logic_vector(to_unsigned( 25, 8)),
9 => std_logic_vector(to_unsigned( 134, 8)),
10 => std_logic_vector(to_unsigned( 31, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 201, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 78, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 43, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 630 then count <= 631; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 228, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 20, 8)),
8 => std_logic_vector(to_unsigned( 32, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 204, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 631 then count <= 632; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 62, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 1, 8)),
11 => std_logic_vector(to_unsigned( 101, 8)),
12 => std_logic_vector(to_unsigned( 215, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 155, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 632 then count <= 633; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 45, 8)),
2 => std_logic_vector(to_unsigned( 64, 8)),
3 => std_logic_vector(to_unsigned( 79, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 87, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 196, 8)),
10 => std_logic_vector(to_unsigned( 215, 8)),
11 => std_logic_vector(to_unsigned( 83, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 59, 8)),
14 => std_logic_vector(to_unsigned( 50, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 633 then count <= 634; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 74, 8)),
4 => std_logic_vector(to_unsigned( 237, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 228, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 221, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 246, 8)),
15 => std_logic_vector(to_unsigned( 32, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 634 then count <= 635; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 156, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 224, 8)),
7 => std_logic_vector(to_unsigned( 164, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 114, 8)),
10 => std_logic_vector(to_unsigned( 35, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 27, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 123, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 635 then count <= 636; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 42, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 254, 8)),
6 => std_logic_vector(to_unsigned( 253, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 40, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 32, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 636 then count <= 637; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 41, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 213, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 216, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 241, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 12, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 637 then count <= 638; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 143, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 40, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 159, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 66, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 243, 8)),
16 => std_logic_vector(to_unsigned( 20, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 638 then count <= 639; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 6, 8)),
3 => std_logic_vector(to_unsigned( 207, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 93, 8)),
6 => std_logic_vector(to_unsigned( 125, 8)),
7 => std_logic_vector(to_unsigned( 14, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 236, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 639 then count <= 640; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 215, 8)),
2 => std_logic_vector(to_unsigned( 228, 8)),
3 => std_logic_vector(to_unsigned( 201, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 74, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 27, 8)),
14 => std_logic_vector(to_unsigned( 126, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 119, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 640 then count <= 641; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 28, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 91, 8)),
6 => std_logic_vector(to_unsigned( 125, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 48, 8)),
9 => std_logic_vector(to_unsigned( 209, 8)),
10 => std_logic_vector(to_unsigned( 162, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 168, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 641 then count <= 642; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 77, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 37, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 118, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 218, 8)),
14 => std_logic_vector(to_unsigned( 119, 8)),
15 => std_logic_vector(to_unsigned( 247, 8)),
16 => std_logic_vector(to_unsigned( 230, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110011
elsif count = 642 then count <= 643; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 45, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 9, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 33, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 22, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 22, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 50, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 643 then count <= 644; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 216, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 228, 8)),
9 => std_logic_vector(to_unsigned( 252, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 226, 8)),
16 => std_logic_vector(to_unsigned( 170, 8)),
17 => std_logic_vector(to_unsigned( 204, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 644 then count <= 645; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 208, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 22, 8)),
8 => std_logic_vector(to_unsigned( 109, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 37, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 209, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 66, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 645 then count <= 646; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 70, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 233, 8)),
6 => std_logic_vector(to_unsigned( 24, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 71, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 646 then count <= 647; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 25, 8)),
5 => std_logic_vector(to_unsigned( 134, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 49, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 1, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 203, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 182, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 647 then count <= 648; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 158, 8)),
2 => std_logic_vector(to_unsigned( 179, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 165, 8)),
5 => std_logic_vector(to_unsigned( 122, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 10, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 219, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 8, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 46, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 648 then count <= 649; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 173, 8)),
12 => std_logic_vector(to_unsigned( 218, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 205, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 649 then count <= 650; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 60, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 10, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 149, 8)),
9 => std_logic_vector(to_unsigned( 41, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 54, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 82, 8)),
15 => std_logic_vector(to_unsigned( 17, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 45, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 650 then count <= 651; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 94, 8)),
2 => std_logic_vector(to_unsigned( 53, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 190, 8)),
11 => std_logic_vector(to_unsigned( 69, 8)),
12 => std_logic_vector(to_unsigned( 180, 8)),
13 => std_logic_vector(to_unsigned( 237, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 651 then count <= 652; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 10, 8)),
3 => std_logic_vector(to_unsigned( 208, 8)),
4 => std_logic_vector(to_unsigned( 6, 8)),
5 => std_logic_vector(to_unsigned( 90, 8)),
6 => std_logic_vector(to_unsigned( 234, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 243, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 16, 8)),
11 => std_logic_vector(to_unsigned( 85, 8)),
12 => std_logic_vector(to_unsigned( 229, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 131, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 652 then count <= 653; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 240, 8)),
3 => std_logic_vector(to_unsigned( 140, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 57, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 98, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 653 then count <= 654; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 20, 8)),
2 => std_logic_vector(to_unsigned( 42, 8)),
3 => std_logic_vector(to_unsigned( 101, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 80, 8)),
7 => std_logic_vector(to_unsigned( 20, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 107, 8)),
11 => std_logic_vector(to_unsigned( 241, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 43, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 218, 8)),
16 => std_logic_vector(to_unsigned( 235, 8)),
17 => std_logic_vector(to_unsigned( 75, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 654 then count <= 655; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 216, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 49, 8)),
4 => std_logic_vector(to_unsigned( 37, 8)),
5 => std_logic_vector(to_unsigned( 227, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 221, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 655 then count <= 656; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 226, 8)),
2 => std_logic_vector(to_unsigned( 249, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 105, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 152, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 156, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 656 then count <= 657; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 116, 8)),
2 => std_logic_vector(to_unsigned( 212, 8)),
3 => std_logic_vector(to_unsigned( 48, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 69, 8)),
9 => std_logic_vector(to_unsigned( 186, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 59, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 136, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 657 then count <= 658; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 152, 8)),
3 => std_logic_vector(to_unsigned( 196, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 150, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 45, 8)),
14 => std_logic_vector(to_unsigned( 232, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 658 then count <= 659; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 2, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 20, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 33, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 659 then count <= 660; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 44, 8)),
2 => std_logic_vector(to_unsigned( 7, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 19, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 82, 8)),
10 => std_logic_vector(to_unsigned( 156, 8)),
11 => std_logic_vector(to_unsigned( 76, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 154, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 167, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 660 then count <= 661; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 210, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 49, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 235, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 51, 8)),
15 => std_logic_vector(to_unsigned( 24, 8)),
16 => std_logic_vector(to_unsigned( 26, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 661 then count <= 662; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 212, 8)),
2 => std_logic_vector(to_unsigned( 197, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 202, 8)),
5 => std_logic_vector(to_unsigned( 221, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 255, 8)),
11 => std_logic_vector(to_unsigned( 221, 8)),
12 => std_logic_vector(to_unsigned( 217, 8)),
13 => std_logic_vector(to_unsigned( 204, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 194, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 222, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 662 then count <= 663; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 236, 8)),
4 => std_logic_vector(to_unsigned( 213, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 44, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 252, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 66, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 42, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110101
elsif count = 663 then count <= 664; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 83, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 229, 8)),
6 => std_logic_vector(to_unsigned( 229, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 24, 8)),
10 => std_logic_vector(to_unsigned( 197, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 74, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 118, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 664 then count <= 665; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 197, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 25, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 159, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 230, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 204, 8)),
15 => std_logic_vector(to_unsigned( 128, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 665 then count <= 666; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 185, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 11, 8)),
8 => std_logic_vector(to_unsigned( 107, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 666 then count <= 667; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 90, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 195, 8)),
8 => std_logic_vector(to_unsigned( 213, 8)),
9 => std_logic_vector(to_unsigned( 245, 8)),
10 => std_logic_vector(to_unsigned( 5, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 79, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 37, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 667 then count <= 668; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 71, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 14, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 14, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 206, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 31, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 210, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 49, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 668 then count <= 669; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 30, 8)),
5 => std_logic_vector(to_unsigned( 156, 8)),
6 => std_logic_vector(to_unsigned( 212, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 189, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 45, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110101
elsif count = 669 then count <= 670; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 252, 8)),
3 => std_logic_vector(to_unsigned( 195, 8)),
4 => std_logic_vector(to_unsigned( 203, 8)),
5 => std_logic_vector(to_unsigned( 215, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 218, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 243, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 1, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 670 then count <= 671; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 170, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 234, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 227, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 227, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 69, 8)),
15 => std_logic_vector(to_unsigned( 99, 8)),
16 => std_logic_vector(to_unsigned( 213, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 211, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 671 then count <= 672; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 85, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 214, 8)),
6 => std_logic_vector(to_unsigned( 219, 8)),
7 => std_logic_vector(to_unsigned( 17, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 107, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 5, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110011
elsif count = 672 then count <= 673; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 170, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 193, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 22, 8)),
10 => std_logic_vector(to_unsigned( 21, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 221, 8)),
13 => std_logic_vector(to_unsigned( 210, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 81, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 673 then count <= 674; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 69, 8)),
2 => std_logic_vector(to_unsigned( 25, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 119, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 228, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 674 then count <= 675; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 186, 8)),
2 => std_logic_vector(to_unsigned( 35, 8)),
3 => std_logic_vector(to_unsigned( 23, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 55, 8)),
6 => std_logic_vector(to_unsigned( 193, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 159, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 50, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 41, 8)),
18 => std_logic_vector(to_unsigned( 149, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 675 then count <= 676; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 10, 8)),
3 => std_logic_vector(to_unsigned( 79, 8)),
4 => std_logic_vector(to_unsigned( 41, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 81, 8)),
7 => std_logic_vector(to_unsigned( 180, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 45, 8)),
10 => std_logic_vector(to_unsigned( 243, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 60, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 36, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 676 then count <= 677; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 158, 8)),
3 => std_logic_vector(to_unsigned( 174, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 12, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 216, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 184, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 218, 8)),
14 => std_logic_vector(to_unsigned( 198, 8)),
15 => std_logic_vector(to_unsigned( 235, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 205, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 677 then count <= 678; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 77, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 102, 8)),
8 => std_logic_vector(to_unsigned( 81, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 77, 8)),
11 => std_logic_vector(to_unsigned( 86, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 179, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 8, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 678 then count <= 679; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 252, 8)),
2 => std_logic_vector(to_unsigned( 20, 8)),
3 => std_logic_vector(to_unsigned( 83, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 231, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 170, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 159, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 197, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 679 then count <= 680; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 146, 8)),
2 => std_logic_vector(to_unsigned( 91, 8)),
3 => std_logic_vector(to_unsigned( 203, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 161, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 198, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 680 then count <= 681; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 127, 8)),
4 => std_logic_vector(to_unsigned( 250, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 31, 8)),
8 => std_logic_vector(to_unsigned( 243, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 242, 8)),
11 => std_logic_vector(to_unsigned( 76, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 219, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 681 then count <= 682; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 125, 8)),
3 => std_logic_vector(to_unsigned( 81, 8)),
4 => std_logic_vector(to_unsigned( 30, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 189, 8)),
7 => std_logic_vector(to_unsigned( 235, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 72, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 175, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110101
elsif count = 682 then count <= 683; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 234, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 58, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 94, 8)),
8 => std_logic_vector(to_unsigned( 130, 8)),
9 => std_logic_vector(to_unsigned( 233, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 20, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 103, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001101
elsif count = 683 then count <= 684; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 166, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 73, 8)),
7 => std_logic_vector(to_unsigned( 84, 8)),
8 => std_logic_vector(to_unsigned( 60, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 229, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 239, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 189, 8)),
15 => std_logic_vector(to_unsigned( 213, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00001111
elsif count = 684 then count <= 685; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 33, 8)),
5 => std_logic_vector(to_unsigned( 142, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 116, 8)),
8 => std_logic_vector(to_unsigned( 135, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 36, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 685 then count <= 686; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 60, 8)),
2 => std_logic_vector(to_unsigned( 32, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 18, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 29, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 33, 8)),
13 => std_logic_vector(to_unsigned( 26, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 40, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 686 then count <= 687; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 118, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 148, 8)),
7 => std_logic_vector(to_unsigned( 60, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 37, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 154, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 687 then count <= 688; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 83, 8)),
2 => std_logic_vector(to_unsigned( 215, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 223, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 56, 8)),
10 => std_logic_vector(to_unsigned( 156, 8)),
11 => std_logic_vector(to_unsigned( 29, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 128, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 688 then count <= 689; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 197, 8)),
2 => std_logic_vector(to_unsigned( 198, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 218, 8)),
7 => std_logic_vector(to_unsigned( 164, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 130, 8)),
10 => std_logic_vector(to_unsigned( 243, 8)),
11 => std_logic_vector(to_unsigned( 150, 8)),
12 => std_logic_vector(to_unsigned( 245, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 249, 8)),
15 => std_logic_vector(to_unsigned( 249, 8)),
16 => std_logic_vector(to_unsigned( 253, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 689 then count <= 690; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 141, 8)),
2 => std_logic_vector(to_unsigned( 176, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 21, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 231, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011010
elsif count = 690 then count <= 691; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 60, 8)),
2 => std_logic_vector(to_unsigned( 31, 8)),
3 => std_logic_vector(to_unsigned( 229, 8)),
4 => std_logic_vector(to_unsigned( 92, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 38, 8)),
8 => std_logic_vector(to_unsigned( 45, 8)),
9 => std_logic_vector(to_unsigned( 26, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 167, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 174, 8)),
17 => std_logic_vector(to_unsigned( 56, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 691 then count <= 692; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 3, 8)),
4 => std_logic_vector(to_unsigned( 214, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 208, 8)),
11 => std_logic_vector(to_unsigned( 65, 8)),
12 => std_logic_vector(to_unsigned( 44, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001101
elsif count = 692 then count <= 693; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 222, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 213, 8)),
5 => std_logic_vector(to_unsigned( 202, 8)),
6 => std_logic_vector(to_unsigned( 127, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 36, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 27, 8)),
12 => std_logic_vector(to_unsigned( 32, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 170, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 693 then count <= 694; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 90, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 84, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 2, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 103, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 694 then count <= 695; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 152, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 163, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 100, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 695 then count <= 696; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 55, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 161, 8)),
8 => std_logic_vector(to_unsigned( 4, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 231, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 237, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 696 then count <= 697; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 30, 8)),
2 => std_logic_vector(to_unsigned( 153, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 1, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 231, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 697 then count <= 698; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 101, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 19, 8)),
10 => std_logic_vector(to_unsigned( 39, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 48, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 1, 8)),
16 => std_logic_vector(to_unsigned( 36, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 698 then count <= 699; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 159, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 108, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 57, 8)),
10 => std_logic_vector(to_unsigned( 87, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 240, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 699 then count <= 700; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 41, 8)),
2 => std_logic_vector(to_unsigned( 96, 8)),
3 => std_logic_vector(to_unsigned( 236, 8)),
4 => std_logic_vector(to_unsigned( 209, 8)),
5 => std_logic_vector(to_unsigned( 146, 8)),
6 => std_logic_vector(to_unsigned( 17, 8)),
7 => std_logic_vector(to_unsigned( 37, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 179, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 28, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 75, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 700 then count <= 701; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 220, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 150, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 14, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 39, 8)),
13 => std_logic_vector(to_unsigned( 222, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 230, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 701 then count <= 702; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 22, 8)),
2 => std_logic_vector(to_unsigned( 194, 8)),
3 => std_logic_vector(to_unsigned( 120, 8)),
4 => std_logic_vector(to_unsigned( 91, 8)),
5 => std_logic_vector(to_unsigned( 253, 8)),
6 => std_logic_vector(to_unsigned( 159, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 233, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 702 then count <= 703; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 59, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 112, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 83, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 107, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 59, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 703 then count <= 704; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 205, 8)),
2 => std_logic_vector(to_unsigned( 218, 8)),
3 => std_logic_vector(to_unsigned( 151, 8)),
4 => std_logic_vector(to_unsigned( 221, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 243, 8)),
7 => std_logic_vector(to_unsigned( 13, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 57, 8)),
12 => std_logic_vector(to_unsigned( 131, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 174, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 704 then count <= 705; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 202, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 193, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 208, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 188, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 209, 8)),
15 => std_logic_vector(to_unsigned( 33, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 187, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 705 then count <= 706; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 159, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 20, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 56, 8)),
9 => std_logic_vector(to_unsigned( 31, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 31, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 235, 8)),
14 => std_logic_vector(to_unsigned( 215, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 706 then count <= 707; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 226, 8)),
2 => std_logic_vector(to_unsigned( 253, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 231, 8)),
10 => std_logic_vector(to_unsigned( 163, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 250, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 707 then count <= 708; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 171, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 238, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 151, 8)),
13 => std_logic_vector(to_unsigned( 221, 8)),
14 => std_logic_vector(to_unsigned( 25, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 708 then count <= 709; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 118, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 36, 8)),
6 => std_logic_vector(to_unsigned( 229, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 151, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 25, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 709 then count <= 710; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 26, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 64, 8)),
5 => std_logic_vector(to_unsigned( 255, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 101, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 209, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 62, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110011
elsif count = 710 then count <= 711; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 84, 8)),
3 => std_logic_vector(to_unsigned( 67, 8)),
4 => std_logic_vector(to_unsigned( 185, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 201, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 39, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 711 then count <= 712; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 155, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 98, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 30, 8)),
9 => std_logic_vector(to_unsigned( 35, 8)),
10 => std_logic_vector(to_unsigned( 54, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 220, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 246, 8)),
16 => std_logic_vector(to_unsigned( 74, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 712 then count <= 713; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 29, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 112, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 52, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 30, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 713 then count <= 714; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 175, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 86, 8)),
6 => std_logic_vector(to_unsigned( 114, 8)),
7 => std_logic_vector(to_unsigned( 41, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 14, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 714 then count <= 715; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 72, 8)),
2 => std_logic_vector(to_unsigned( 54, 8)),
3 => std_logic_vector(to_unsigned( 156, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 3, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 163, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 33, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 715 then count <= 716; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 101, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 236, 8)),
8 => std_logic_vector(to_unsigned( 61, 8)),
9 => std_logic_vector(to_unsigned( 111, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 54, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 255, 8)),
14 => std_logic_vector(to_unsigned( 34, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 54, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 716 then count <= 717; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 212, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 36, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 164, 8)),
8 => std_logic_vector(to_unsigned( 153, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 219, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 8, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 717 then count <= 718; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 66, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 103, 8)),
6 => std_logic_vector(to_unsigned( 160, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 204, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 29, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 55, 8)),
14 => std_logic_vector(to_unsigned( 208, 8)),
15 => std_logic_vector(to_unsigned( 33, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 718 then count <= 719; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 160, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 184, 8)),
5 => std_logic_vector(to_unsigned( 10, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 166, 8)),
9 => std_logic_vector(to_unsigned( 199, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 40, 8)),
12 => std_logic_vector(to_unsigned( 42, 8)),
13 => std_logic_vector(to_unsigned( 207, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 170, 8)),
16 => std_logic_vector(to_unsigned( 238, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 719 then count <= 720; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 67, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 17, 8)),
4 => std_logic_vector(to_unsigned( 79, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 21, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 193, 8)),
9 => std_logic_vector(to_unsigned( 9, 8)),
10 => std_logic_vector(to_unsigned( 71, 8)),
11 => std_logic_vector(to_unsigned( 30, 8)),
12 => std_logic_vector(to_unsigned( 48, 8)),
13 => std_logic_vector(to_unsigned( 47, 8)),
14 => std_logic_vector(to_unsigned( 31, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 75, 8)),
18 => std_logic_vector(to_unsigned( 70, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 720 then count <= 721; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 220, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 217, 8)),
5 => std_logic_vector(to_unsigned( 4, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 237, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 173, 8)),
12 => std_logic_vector(to_unsigned( 88, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 206, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 721 then count <= 722; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 45, 8)),
2 => std_logic_vector(to_unsigned( 241, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 231, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 184, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 222, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 131, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 722 then count <= 723; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 49, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 60, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 14, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 112, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 157, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 66, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 723 then count <= 724; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 44, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 32, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 254, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 55, 8)),
9 => std_logic_vector(to_unsigned( 206, 8)),
10 => std_logic_vector(to_unsigned( 254, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 66, 8)),
14 => std_logic_vector(to_unsigned( 3, 8)),
15 => std_logic_vector(to_unsigned( 25, 8)),
16 => std_logic_vector(to_unsigned( 47, 8)),
17 => std_logic_vector(to_unsigned( 41, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 724 then count <= 725; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 8, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 165, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 206, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 235, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 218, 8)),
15 => std_logic_vector(to_unsigned( 234, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 725 then count <= 726; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 3, 8)),
3 => std_logic_vector(to_unsigned( 171, 8)),
4 => std_logic_vector(to_unsigned( 28, 8)),
5 => std_logic_vector(to_unsigned( 198, 8)),
6 => std_logic_vector(to_unsigned( 2, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 29, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 28, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 23, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 232, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 36, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 726 then count <= 727; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 162, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 220, 8)),
7 => std_logic_vector(to_unsigned( 208, 8)),
8 => std_logic_vector(to_unsigned( 8, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 36, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 170, 8)),
16 => std_logic_vector(to_unsigned( 105, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 727 then count <= 728; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 190, 8)),
2 => std_logic_vector(to_unsigned( 48, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 119, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 10, 8)),
8 => std_logic_vector(to_unsigned( 59, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 77, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 5, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 728 then count <= 729; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 139, 8)),
2 => std_logic_vector(to_unsigned( 244, 8)),
3 => std_logic_vector(to_unsigned( 208, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 10, 8)),
6 => std_logic_vector(to_unsigned( 22, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 32, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 163, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 158, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 200, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110000
elsif count = 729 then count <= 730; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 94, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 88, 8)),
7 => std_logic_vector(to_unsigned( 48, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 41, 8)),
10 => std_logic_vector(to_unsigned( 243, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 58, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 7, 8)),
16 => std_logic_vector(to_unsigned( 47, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101110
elsif count = 730 then count <= 731; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 244, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 38, 8)),
6 => std_logic_vector(to_unsigned( 235, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 201, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 205, 8)),
11 => std_logic_vector(to_unsigned( 247, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 45, 8)),
14 => std_logic_vector(to_unsigned( 18, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 207, 8)),
17 => std_logic_vector(to_unsigned( 52, 8)),
18 => std_logic_vector(to_unsigned( 198, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 731 then count <= 732; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 239, 8)),
2 => std_logic_vector(to_unsigned( 235, 8)),
3 => std_logic_vector(to_unsigned( 37, 8)),
4 => std_logic_vector(to_unsigned( 165, 8)),
5 => std_logic_vector(to_unsigned( 100, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 56, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 111, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 24, 8)),
14 => std_logic_vector(to_unsigned( 186, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 732 then count <= 733; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 158, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 182, 8)),
7 => std_logic_vector(to_unsigned( 154, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 126, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 70, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 39, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 733 then count <= 734; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 146, 8)),
2 => std_logic_vector(to_unsigned( 228, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 13, 8)),
11 => std_logic_vector(to_unsigned( 13, 8)),
12 => std_logic_vector(to_unsigned( 57, 8)),
13 => std_logic_vector(to_unsigned( 6, 8)),
14 => std_logic_vector(to_unsigned( 62, 8)),
15 => std_logic_vector(to_unsigned( 143, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001110
elsif count = 734 then count <= 735; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 198, 8)),
2 => std_logic_vector(to_unsigned( 142, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 61, 8)),
5 => std_logic_vector(to_unsigned( 7, 8)),
6 => std_logic_vector(to_unsigned( 232, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 156, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 247, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 735 then count <= 736; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 238, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 67, 8)),
4 => std_logic_vector(to_unsigned( 56, 8)),
5 => std_logic_vector(to_unsigned( 204, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 173, 8)),
14 => std_logic_vector(to_unsigned( 100, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 41, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 736 then count <= 737; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 109, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 132, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 251, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 41, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 737 then count <= 738; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 247, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 241, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 11, 8)),
6 => std_logic_vector(to_unsigned( 10, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 231, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 238, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 738 then count <= 739; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 218, 8)),
3 => std_logic_vector(to_unsigned( 200, 8)),
4 => std_logic_vector(to_unsigned( 118, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 209, 8)),
7 => std_logic_vector(to_unsigned( 204, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 205, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 61, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 212, 8)),
16 => std_logic_vector(to_unsigned( 15, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 739 then count <= 740; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 146, 8)),
2 => std_logic_vector(to_unsigned( 34, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 73, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 123, 8)),
7 => std_logic_vector(to_unsigned( 238, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 116, 8)),
11 => std_logic_vector(to_unsigned( 4, 8)),
12 => std_logic_vector(to_unsigned( 246, 8)),
13 => std_logic_vector(to_unsigned( 219, 8)),
14 => std_logic_vector(to_unsigned( 100, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 33, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 740 then count <= 741; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 227, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 214, 8)),
5 => std_logic_vector(to_unsigned( 59, 8)),
6 => std_logic_vector(to_unsigned( 159, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 109, 8)),
9 => std_logic_vector(to_unsigned( 225, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 183, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 134, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 741 then count <= 742; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 3, 8)),
4 => std_logic_vector(to_unsigned( 43, 8)),
5 => std_logic_vector(to_unsigned( 119, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 219, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 222, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 181, 8)),
15 => std_logic_vector(to_unsigned( 35, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 742 then count <= 743; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 117, 8)),
6 => std_logic_vector(to_unsigned( 62, 8)),
7 => std_logic_vector(to_unsigned( 98, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 72, 8)),
10 => std_logic_vector(to_unsigned( 221, 8)),
11 => std_logic_vector(to_unsigned( 120, 8)),
12 => std_logic_vector(to_unsigned( 59, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 224, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 743 then count <= 744; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 254, 8)),
2 => std_logic_vector(to_unsigned( 2, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 59, 8)),
11 => std_logic_vector(to_unsigned( 218, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 194, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 193, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 744 then count <= 745; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 217, 8)),
2 => std_logic_vector(to_unsigned( 5, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 9, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 45, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 166, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 183, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 745 then count <= 746; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 146, 8)),
2 => std_logic_vector(to_unsigned( 219, 8)),
3 => std_logic_vector(to_unsigned( 157, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 217, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100100
elsif count = 746 then count <= 747; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 44, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 129, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 178, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 747 then count <= 748; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 64, 8)),
5 => std_logic_vector(to_unsigned( 215, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 249, 8)),
11 => std_logic_vector(to_unsigned( 208, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 748 then count <= 749; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 227, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 1, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 112, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 42, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 98, 8)),
13 => std_logic_vector(to_unsigned( 141, 8)),
14 => std_logic_vector(to_unsigned( 128, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 749 then count <= 750; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 214, 8)),
4 => std_logic_vector(to_unsigned( 226, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 231, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 246, 8)),
10 => std_logic_vector(to_unsigned( 45, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 230, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 750 then count <= 751; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 170, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 220, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 182, 8)),
10 => std_logic_vector(to_unsigned( 245, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 156, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 170, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 106, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 751 then count <= 752; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 9, 8)),
3 => std_logic_vector(to_unsigned( 46, 8)),
4 => std_logic_vector(to_unsigned( 209, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 249, 8)),
7 => std_logic_vector(to_unsigned( 56, 8)),
8 => std_logic_vector(to_unsigned( 241, 8)),
9 => std_logic_vector(to_unsigned( 77, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 59, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 196, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 220, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 752 then count <= 753; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 100, 8)),
6 => std_logic_vector(to_unsigned( 95, 8)),
7 => std_logic_vector(to_unsigned( 230, 8)),
8 => std_logic_vector(to_unsigned( 252, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 239, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 191, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 753 then count <= 754; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 119, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 18, 8)),
8 => std_logic_vector(to_unsigned( 227, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 217, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 173, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 172, 8)),
16 => std_logic_vector(to_unsigned( 153, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 754 then count <= 755; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 221, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 189, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 101, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 4, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 18, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 210, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 755 then count <= 756; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 40, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 208, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 179, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 756 then count <= 757; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 221, 8)),
3 => std_logic_vector(to_unsigned( 178, 8)),
4 => std_logic_vector(to_unsigned( 45, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 156, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 66, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 163, 8)),
12 => std_logic_vector(to_unsigned( 52, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 757 then count <= 758; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 129, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 60, 8)),
9 => std_logic_vector(to_unsigned( 138, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 185, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 758 then count <= 759; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 206, 8)),
2 => std_logic_vector(to_unsigned( 215, 8)),
3 => std_logic_vector(to_unsigned( 83, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 220, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 3, 8)),
8 => std_logic_vector(to_unsigned( 28, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 236, 8)),
12 => std_logic_vector(to_unsigned( 12, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 180, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 759 then count <= 760; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 187, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 124, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 164, 8)),
9 => std_logic_vector(to_unsigned( 213, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 181, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 231, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 760 then count <= 761; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 205, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 27, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 80, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 3, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 761 then count <= 762; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 129, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 110, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 173, 8)),
12 => std_logic_vector(to_unsigned( 151, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 236, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 246, 8)),
17 => std_logic_vector(to_unsigned( 118, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 762 then count <= 763; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 30, 8)),
4 => std_logic_vector(to_unsigned( 7, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 141, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 763 then count <= 764; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 249, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 32, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 94, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 141, 8)),
15 => std_logic_vector(to_unsigned( 215, 8)),
16 => std_logic_vector(to_unsigned( 131, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 764 then count <= 765; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 16, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 55, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 22, 8)),
7 => std_logic_vector(to_unsigned( 195, 8)),
8 => std_logic_vector(to_unsigned( 120, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 47, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 176, 8)),
14 => std_logic_vector(to_unsigned( 238, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 765 then count <= 766; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 4, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 41, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 112, 8)),
11 => std_logic_vector(to_unsigned( 249, 8)),
12 => std_logic_vector(to_unsigned( 230, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001100
elsif count = 766 then count <= 767; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 216, 8)),
2 => std_logic_vector(to_unsigned( 192, 8)),
3 => std_logic_vector(to_unsigned( 41, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 164, 8)),
6 => std_logic_vector(to_unsigned( 71, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 21, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 38, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 18, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 767 then count <= 768; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 76, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 36, 8)),
6 => std_logic_vector(to_unsigned( 1, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 34, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 95, 8)),
14 => std_logic_vector(to_unsigned( 211, 8)),
15 => std_logic_vector(to_unsigned( 81, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100010
elsif count = 768 then count <= 769; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 56, 8)),
4 => std_logic_vector(to_unsigned( 184, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 245, 8)),
7 => std_logic_vector(to_unsigned( 211, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 21, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 145, 8)),
17 => std_logic_vector(to_unsigned( 49, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 769 then count <= 770; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 76, 8)),
4 => std_logic_vector(to_unsigned( 90, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 210, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 149, 8)),
9 => std_logic_vector(to_unsigned( 182, 8)),
10 => std_logic_vector(to_unsigned( 179, 8)),
11 => std_logic_vector(to_unsigned( 3, 8)),
12 => std_logic_vector(to_unsigned( 57, 8)),
13 => std_logic_vector(to_unsigned( 43, 8)),
14 => std_logic_vector(to_unsigned( 222, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 770 then count <= 771; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 99, 8)),
2 => std_logic_vector(to_unsigned( 51, 8)),
3 => std_logic_vector(to_unsigned( 178, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 249, 8)),
7 => std_logic_vector(to_unsigned( 181, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 198, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 17, 8)),
14 => std_logic_vector(to_unsigned( 47, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 771 then count <= 772; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 229, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 8, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 173, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 74, 8)),
14 => std_logic_vector(to_unsigned( 67, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 119, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100010
elsif count = 772 then count <= 773; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 226, 8)),
6 => std_logic_vector(to_unsigned( 73, 8)),
7 => std_logic_vector(to_unsigned( 236, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 240, 8)),
10 => std_logic_vector(to_unsigned( 115, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 198, 8)),
13 => std_logic_vector(to_unsigned( 34, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 220, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 773 then count <= 774; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 174, 8)),
8 => std_logic_vector(to_unsigned( 85, 8)),
9 => std_logic_vector(to_unsigned( 5, 8)),
10 => std_logic_vector(to_unsigned( 124, 8)),
11 => std_logic_vector(to_unsigned( 107, 8)),
12 => std_logic_vector(to_unsigned( 154, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 246, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 774 then count <= 775; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 177, 8)),
8 => std_logic_vector(to_unsigned( 91, 8)),
9 => std_logic_vector(to_unsigned( 137, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 216, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 97, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 775 then count <= 776; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 47, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 234, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 142, 8)),
7 => std_logic_vector(to_unsigned( 16, 8)),
8 => std_logic_vector(to_unsigned( 52, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 68, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 9, 8)),
14 => std_logic_vector(to_unsigned( 3, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110110
elsif count = 776 then count <= 777; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 171, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 25, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 204, 8)),
10 => std_logic_vector(to_unsigned( 122, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 116, 8)),
13 => std_logic_vector(to_unsigned( 98, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 136, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110101
elsif count = 777 then count <= 778; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 212, 8)),
2 => std_logic_vector(to_unsigned( 251, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 25, 8)),
5 => std_logic_vector(to_unsigned( 88, 8)),
6 => std_logic_vector(to_unsigned( 238, 8)),
7 => std_logic_vector(to_unsigned( 103, 8)),
8 => std_logic_vector(to_unsigned( 171, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 40, 8)),
13 => std_logic_vector(to_unsigned( 79, 8)),
14 => std_logic_vector(to_unsigned( 165, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 778 then count <= 779; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 207, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 39, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 66, 8)),
8 => std_logic_vector(to_unsigned( 234, 8)),
9 => std_logic_vector(to_unsigned( 148, 8)),
10 => std_logic_vector(to_unsigned( 169, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 10, 8)),
13 => std_logic_vector(to_unsigned( 210, 8)),
14 => std_logic_vector(to_unsigned( 45, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 222, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 779 then count <= 780; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 248, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 104, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 177, 8)),
8 => std_logic_vector(to_unsigned( 52, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 54, 8)),
11 => std_logic_vector(to_unsigned( 33, 8)),
12 => std_logic_vector(to_unsigned( 5, 8)),
13 => std_logic_vector(to_unsigned( 15, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 25, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 48, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 780 then count <= 781; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 211, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 28, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 31, 8)),
7 => std_logic_vector(to_unsigned( 247, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 224, 8)),
10 => std_logic_vector(to_unsigned( 210, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 238, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 141, 8)),
17 => std_logic_vector(to_unsigned( 181, 8)),
18 => std_logic_vector(to_unsigned( 185, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 781 then count <= 782; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 21, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 13, 8)),
11 => std_logic_vector(to_unsigned( 221, 8)),
12 => std_logic_vector(to_unsigned( 220, 8)),
13 => std_logic_vector(to_unsigned( 50, 8)),
14 => std_logic_vector(to_unsigned( 82, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 77, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 128, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 782 then count <= 783; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 17, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 31, 8)),
7 => std_logic_vector(to_unsigned( 38, 8)),
8 => std_logic_vector(to_unsigned( 3, 8)),
9 => std_logic_vector(to_unsigned( 21, 8)),
10 => std_logic_vector(to_unsigned( 16, 8)),
11 => std_logic_vector(to_unsigned( 36, 8)),
12 => std_logic_vector(to_unsigned( 1, 8)),
13 => std_logic_vector(to_unsigned( 179, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 227, 8)),
16 => std_logic_vector(to_unsigned( 248, 8)),
17 => std_logic_vector(to_unsigned( 36, 8)),
18 => std_logic_vector(to_unsigned( 34, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 783 then count <= 784; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 223, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 75, 8)),
5 => std_logic_vector(to_unsigned( 228, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 116, 8)),
11 => std_logic_vector(to_unsigned( 2, 8)),
12 => std_logic_vector(to_unsigned( 96, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 182, 8)),
16 => std_logic_vector(to_unsigned( 73, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 784 then count <= 785; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 224, 8)),
2 => std_logic_vector(to_unsigned( 32, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 184, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 4, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 63, 8)),
13 => std_logic_vector(to_unsigned( 178, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 185, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001100
elsif count = 785 then count <= 786; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 185, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 23, 8)),
5 => std_logic_vector(to_unsigned( 180, 8)),
6 => std_logic_vector(to_unsigned( 15, 8)),
7 => std_logic_vector(to_unsigned( 154, 8)),
8 => std_logic_vector(to_unsigned( 127, 8)),
9 => std_logic_vector(to_unsigned( 213, 8)),
10 => std_logic_vector(to_unsigned( 22, 8)),
11 => std_logic_vector(to_unsigned( 176, 8)),
12 => std_logic_vector(to_unsigned( 51, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 6, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 35, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 786 then count <= 787; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 131, 8)),
4 => std_logic_vector(to_unsigned( 2, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 28, 8)),
7 => std_logic_vector(to_unsigned( 50, 8)),
8 => std_logic_vector(to_unsigned( 255, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 31, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 21, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 3, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 787 then count <= 788; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 204, 8)),
4 => std_logic_vector(to_unsigned( 181, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 112, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 52, 8)),
15 => std_logic_vector(to_unsigned( 167, 8)),
16 => std_logic_vector(to_unsigned( 225, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 788 then count <= 789; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 249, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 204, 8)),
6 => std_logic_vector(to_unsigned( 148, 8)),
7 => std_logic_vector(to_unsigned( 245, 8)),
8 => std_logic_vector(to_unsigned( 189, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 129, 8)),
12 => std_logic_vector(to_unsigned( 232, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 236, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 24, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 193, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 789 then count <= 790; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 37, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 222, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 55, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 255, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 58, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 790 then count <= 791; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 71, 8)),
3 => std_logic_vector(to_unsigned( 199, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 238, 8)),
7 => std_logic_vector(to_unsigned( 254, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 86, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 175, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 8, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 791 then count <= 792; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 55, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 234, 8)),
5 => std_logic_vector(to_unsigned( 122, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 17, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 232, 8)),
11 => std_logic_vector(to_unsigned( 167, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 218, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 121, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 792 then count <= 793; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 17, 8)),
2 => std_logic_vector(to_unsigned( 192, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 59, 8)),
5 => std_logic_vector(to_unsigned( 203, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 233, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 229, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 190, 8)),
14 => std_logic_vector(to_unsigned( 21, 8)),
15 => std_logic_vector(to_unsigned( 232, 8)),
16 => std_logic_vector(to_unsigned( 63, 8)),
17 => std_logic_vector(to_unsigned( 190, 8)),
18 => std_logic_vector(to_unsigned( 70, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 793 then count <= 794; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 211, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 41, 8)),
6 => std_logic_vector(to_unsigned( 79, 8)),
7 => std_logic_vector(to_unsigned( 83, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 43, 8)),
12 => std_logic_vector(to_unsigned( 0, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 794 then count <= 795; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 152, 8)),
3 => std_logic_vector(to_unsigned( 89, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 159, 8)),
9 => std_logic_vector(to_unsigned( 191, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 27, 8)),
12 => std_logic_vector(to_unsigned( 203, 8)),
13 => std_logic_vector(to_unsigned( 173, 8)),
14 => std_logic_vector(to_unsigned( 26, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 246, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 795 then count <= 796; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 69, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 39, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 13, 8)),
8 => std_logic_vector(to_unsigned( 27, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 72, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 43, 8)),
14 => std_logic_vector(to_unsigned( 188, 8)),
15 => std_logic_vector(to_unsigned( 215, 8)),
16 => std_logic_vector(to_unsigned( 239, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 796 then count <= 797; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 33, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 33, 8)),
8 => std_logic_vector(to_unsigned( 8, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 189, 8)),
11 => std_logic_vector(to_unsigned( 24, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 194, 8)),
15 => std_logic_vector(to_unsigned( 30, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 59, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 797 then count <= 798; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 85, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 247, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 237, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 241, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 69, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 250, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 52, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 218, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 798 then count <= 799; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 51, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 60, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 28, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 61, 8)),
16 => std_logic_vector(to_unsigned( 46, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 799 then count <= 800; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 240, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 208, 8)),
5 => std_logic_vector(to_unsigned( 231, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 246, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 800 then count <= 801; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 255, 8)),
2 => std_logic_vector(to_unsigned( 200, 8)),
3 => std_logic_vector(to_unsigned( 197, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 188, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 165, 8)),
15 => std_logic_vector(to_unsigned( 12, 8)),
16 => std_logic_vector(to_unsigned( 244, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 801 then count <= 802; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 255, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 224, 8)),
13 => std_logic_vector(to_unsigned( 173, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 218, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 802 then count <= 803; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 206, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 110, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 214, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 152, 8)),
13 => std_logic_vector(to_unsigned( 223, 8)),
14 => std_logic_vector(to_unsigned( 255, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 803 then count <= 804; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 193, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 49, 8)),
9 => std_logic_vector(to_unsigned( 110, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 17, 8)),
12 => std_logic_vector(to_unsigned( 242, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 250, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 196, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 206, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010101
elsif count = 804 then count <= 805; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 109, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 133, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 247, 8)),
11 => std_logic_vector(to_unsigned( 216, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 24, 8)),
14 => std_logic_vector(to_unsigned( 56, 8)),
15 => std_logic_vector(to_unsigned( 23, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 62, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 805 then count <= 806; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 72, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 43, 8)),
5 => std_logic_vector(to_unsigned( 2, 8)),
6 => std_logic_vector(to_unsigned( 21, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 59, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 132, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 806 then count <= 807; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 41, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 3, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 10, 8)),
7 => std_logic_vector(to_unsigned( 77, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 18, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 131, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 807 then count <= 808; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 220, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 76, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 67, 8)),
8 => std_logic_vector(to_unsigned( 182, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 210, 8)),
13 => std_logic_vector(to_unsigned( 28, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 206, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 808 then count <= 809; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 215, 8)),
3 => std_logic_vector(to_unsigned( 193, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 158, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 215, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 253, 8)),
10 => std_logic_vector(to_unsigned( 228, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 204, 8)),
14 => std_logic_vector(to_unsigned( 57, 8)),
15 => std_logic_vector(to_unsigned( 10, 8)),
16 => std_logic_vector(to_unsigned( 17, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 809 then count <= 810; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 40, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 68, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 232, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 229, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 42, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 231, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 810 then count <= 811; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 108, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 7, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 54, 8)),
9 => std_logic_vector(to_unsigned( 57, 8)),
10 => std_logic_vector(to_unsigned( 230, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 13, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 2, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 74, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001011
elsif count = 811 then count <= 812; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 181, 8)),
9 => std_logic_vector(to_unsigned( 137, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 181, 8)),
12 => std_logic_vector(to_unsigned( 33, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 62, 8)),
15 => std_logic_vector(to_unsigned( 234, 8)),
16 => std_logic_vector(to_unsigned( 249, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 812 then count <= 813; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 162, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 217, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 211, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 42, 8)),
10 => std_logic_vector(to_unsigned( 63, 8)),
11 => std_logic_vector(to_unsigned( 203, 8)),
12 => std_logic_vector(to_unsigned( 157, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 196, 8)),
17 => std_logic_vector(to_unsigned( 197, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 813 then count <= 814; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 219, 8)),
3 => std_logic_vector(to_unsigned( 237, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 16, 8)),
6 => std_logic_vector(to_unsigned( 24, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 132, 8)),
9 => std_logic_vector(to_unsigned( 226, 8)),
10 => std_logic_vector(to_unsigned( 112, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 81, 8)),
16 => std_logic_vector(to_unsigned( 196, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 814 then count <= 815; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 32, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 16, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 9, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 228, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 15, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 92, 8)),
12 => std_logic_vector(to_unsigned( 237, 8)),
13 => std_logic_vector(to_unsigned( 204, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 232, 8)),
17 => std_logic_vector(to_unsigned( 33, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00010111
elsif count = 815 then count <= 816; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 240, 8)),
2 => std_logic_vector(to_unsigned( 206, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 220, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 77, 8)),
13 => std_logic_vector(to_unsigned( 141, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 248, 8)),
16 => std_logic_vector(to_unsigned( 174, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 816 then count <= 817; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 133, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 203, 8)),
11 => std_logic_vector(to_unsigned( 181, 8)),
12 => std_logic_vector(to_unsigned( 77, 8)),
13 => std_logic_vector(to_unsigned( 14, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001110
elsif count = 817 then count <= 818; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 193, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 164, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 170, 8)),
9 => std_logic_vector(to_unsigned( 141, 8)),
10 => std_logic_vector(to_unsigned( 47, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 204, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 189, 8)),
18 => std_logic_vector(to_unsigned( 198, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 818 then count <= 819; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 39, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 49, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 99, 8)),
10 => std_logic_vector(to_unsigned( 206, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 210, 8)),
13 => std_logic_vector(to_unsigned( 47, 8)),
14 => std_logic_vector(to_unsigned( 57, 8)),
15 => std_logic_vector(to_unsigned( 193, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 819 then count <= 820; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 92, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 80, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 190, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 207, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 184, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 218, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 820 then count <= 821; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 224, 8)),
2 => std_logic_vector(to_unsigned( 21, 8)),
3 => std_logic_vector(to_unsigned( 56, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 181, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 164, 8)),
8 => std_logic_vector(to_unsigned( 220, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 200, 8)),
12 => std_logic_vector(to_unsigned( 42, 8)),
13 => std_logic_vector(to_unsigned( 4, 8)),
14 => std_logic_vector(to_unsigned( 228, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 821 then count <= 822; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 145, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 202, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 82, 8)),
9 => std_logic_vector(to_unsigned( 84, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 233, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 33, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 822 then count <= 823; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 45, 8)),
3 => std_logic_vector(to_unsigned( 86, 8)),
4 => std_logic_vector(to_unsigned( 164, 8)),
5 => std_logic_vector(to_unsigned( 164, 8)),
6 => std_logic_vector(to_unsigned( 216, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 89, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 79, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 199, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 823 then count <= 824; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 207, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 18, 8)),
6 => std_logic_vector(to_unsigned( 211, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 241, 8)),
9 => std_logic_vector(to_unsigned( 254, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 229, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 234, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 824 then count <= 825; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 223, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 23, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 255, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 74, 8)),
13 => std_logic_vector(to_unsigned( 95, 8)),
14 => std_logic_vector(to_unsigned( 146, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 232, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 825 then count <= 826; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 220, 8)),
2 => std_logic_vector(to_unsigned( 63, 8)),
3 => std_logic_vector(to_unsigned( 243, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 134, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 195, 8)),
8 => std_logic_vector(to_unsigned( 253, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 37, 8)),
14 => std_logic_vector(to_unsigned( 228, 8)),
15 => std_logic_vector(to_unsigned( 242, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010011
elsif count = 826 then count <= 827; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 10, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 134, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 168, 8)),
8 => std_logic_vector(to_unsigned( 132, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 66, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 123, 8)),
18 => std_logic_vector(to_unsigned( 46, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 827 then count <= 828; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 0, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 215, 8)),
5 => std_logic_vector(to_unsigned( 78, 8)),
6 => std_logic_vector(to_unsigned( 194, 8)),
7 => std_logic_vector(to_unsigned( 250, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 156, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 193, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 828 then count <= 829; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 215, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 133, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 54, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 220, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 147, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 829 then count <= 830; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 31, 8)),
2 => std_logic_vector(to_unsigned( 212, 8)),
3 => std_logic_vector(to_unsigned( 14, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 233, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 39, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 239, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 229, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 830 then count <= 831; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 36, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 139, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 47, 8)),
16 => std_logic_vector(to_unsigned( 177, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 831 then count <= 832; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 16, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 116, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 72, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 249, 8)),
12 => std_logic_vector(to_unsigned( 109, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 46, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 832 then count <= 833; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 165, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 88, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 65, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 46, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 24, 8)),
14 => std_logic_vector(to_unsigned( 21, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 833 then count <= 834; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 213, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 244, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 208, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 70, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 195, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 834 then count <= 835; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 211, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 19, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 234, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 190, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 30, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 21, 8)),
17 => std_logic_vector(to_unsigned( 207, 8)),
18 => std_logic_vector(to_unsigned( 38, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 835 then count <= 836; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 188, 8)),
3 => std_logic_vector(to_unsigned( 5, 8)),
4 => std_logic_vector(to_unsigned( 235, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 239, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 232, 8)),
10 => std_logic_vector(to_unsigned( 200, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 211, 8)),
13 => std_logic_vector(to_unsigned( 229, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 240, 8)),
16 => std_logic_vector(to_unsigned( 206, 8)),
17 => std_logic_vector(to_unsigned( 211, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 836 then count <= 837; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 20, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 151, 8)),
9 => std_logic_vector(to_unsigned( 23, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 60, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 74, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 54, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 837 then count <= 838; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 187, 8)),
5 => std_logic_vector(to_unsigned( 233, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 191, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 136, 8)),
11 => std_logic_vector(to_unsigned( 27, 8)),
12 => std_logic_vector(to_unsigned( 110, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 163, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 838 then count <= 839; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 201, 8)),
4 => std_logic_vector(to_unsigned( 49, 8)),
5 => std_logic_vector(to_unsigned( 249, 8)),
6 => std_logic_vector(to_unsigned( 16, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 200, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 183, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 196, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 839 then count <= 840; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 227, 8)),
2 => std_logic_vector(to_unsigned( 194, 8)),
3 => std_logic_vector(to_unsigned( 112, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 217, 8)),
6 => std_logic_vector(to_unsigned( 123, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 179, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 228, 8)),
11 => std_logic_vector(to_unsigned( 33, 8)),
12 => std_logic_vector(to_unsigned( 34, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 840 then count <= 841; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 98, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 841 then count <= 842; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 38, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 227, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 248, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 14, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 842 then count <= 843; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 231, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 207, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 195, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 198, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 217, 8)),
17 => std_logic_vector(to_unsigned( 208, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 843 then count <= 844; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 23, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 163, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 2, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 23, 8)),
10 => std_logic_vector(to_unsigned( 212, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 74, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 844 then count <= 845; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 190, 8)),
3 => std_logic_vector(to_unsigned( 39, 8)),
4 => std_logic_vector(to_unsigned( 249, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 62, 8)),
12 => std_logic_vector(to_unsigned( 33, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 845 then count <= 846; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 66, 8)),
2 => std_logic_vector(to_unsigned( 192, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 245, 8)),
5 => std_logic_vector(to_unsigned( 241, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 249, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 101, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 151, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 78, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 846 then count <= 847; RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 221, 8)),
3 => std_logic_vector(to_unsigned( 216, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 241, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 242, 8)),
11 => std_logic_vector(to_unsigned( 245, 8)),
12 => std_logic_vector(to_unsigned( 249, 8)),
13 => std_logic_vector(to_unsigned( 150, 8)),
14 => std_logic_vector(to_unsigned( 238, 8)),
15 => std_logic_vector(to_unsigned( 136, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 214, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 847 then count <= 848; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 69, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 253, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 91, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 56, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 61, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 229, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 91, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 848 then count <= 849; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 185, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 195, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 211, 8)),
7 => std_logic_vector(to_unsigned( 60, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 225, 8)),
10 => std_logic_vector(to_unsigned( 136, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 50, 8)),
13 => std_logic_vector(to_unsigned( 173, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 204, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 849 then count <= 850; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 1, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 240, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 49, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 850 then count <= 851; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 130, 8)),
2 => std_logic_vector(to_unsigned( 219, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 245, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 216, 8)),
8 => std_logic_vector(to_unsigned( 106, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 240, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 152, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 190, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 851 then count <= 852; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 226, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 184, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 209, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 150, 8)),
14 => std_logic_vector(to_unsigned( 34, 8)),
15 => std_logic_vector(to_unsigned( 209, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 60, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 852 then count <= 853; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 163, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 8, 8)),
9 => std_logic_vector(to_unsigned( 177, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 128, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 98, 8)),
17 => std_logic_vector(to_unsigned( 200, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110110
elsif count = 853 then count <= 854; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 174, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 183, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 37, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 243, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 102, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 854 then count <= 855; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 141, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 193, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 243, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 30, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 216, 8)),
13 => std_logic_vector(to_unsigned( 4, 8)),
14 => std_logic_vector(to_unsigned( 204, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 855 then count <= 856; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 80, 8)),
2 => std_logic_vector(to_unsigned( 55, 8)),
3 => std_logic_vector(to_unsigned( 8, 8)),
4 => std_logic_vector(to_unsigned( 64, 8)),
5 => std_logic_vector(to_unsigned( 82, 8)),
6 => std_logic_vector(to_unsigned( 53, 8)),
7 => std_logic_vector(to_unsigned( 223, 8)),
8 => std_logic_vector(to_unsigned( 249, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 64, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 121, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 856 then count <= 857; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 43, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 86, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 151, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 44, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 130, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 857 then count <= 858; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 62, 8)),
3 => std_logic_vector(to_unsigned( 254, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 63, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 10, 8)),
10 => std_logic_vector(to_unsigned( 0, 8)),
11 => std_logic_vector(to_unsigned( 199, 8)),
12 => std_logic_vector(to_unsigned( 222, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 159, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 858 then count <= 859; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 205, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 112, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 56, 8)),
12 => std_logic_vector(to_unsigned( 10, 8)),
13 => std_logic_vector(to_unsigned( 195, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 164, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011001
elsif count = 859 then count <= 860; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 24, 8)),
10 => std_logic_vector(to_unsigned( 232, 8)),
11 => std_logic_vector(to_unsigned( 87, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 56, 8)),
15 => std_logic_vector(to_unsigned( 225, 8)),
16 => std_logic_vector(to_unsigned( 213, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 860 then count <= 861; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 158, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 245, 8)),
16 => std_logic_vector(to_unsigned( 241, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 861 then count <= 862; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 242, 8)),
3 => std_logic_vector(to_unsigned( 205, 8)),
4 => std_logic_vector(to_unsigned( 29, 8)),
5 => std_logic_vector(to_unsigned( 170, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 53, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 43, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 80, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 862 then count <= 863; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 156, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 98, 8)),
8 => std_logic_vector(to_unsigned( 41, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 16, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 182, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 863 then count <= 864; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 197, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 116, 8)),
5 => std_logic_vector(to_unsigned( 14, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 15, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 248, 8)),
14 => std_logic_vector(to_unsigned( 77, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 864 then count <= 865; RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 155, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 58, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 53, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 29, 8)),
12 => std_logic_vector(to_unsigned( 245, 8)),
13 => std_logic_vector(to_unsigned( 209, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 40, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 865 then count <= 866; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 45, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 177, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 27, 8)),
14 => std_logic_vector(to_unsigned( 63, 8)),
15 => std_logic_vector(to_unsigned( 35, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 866 then count <= 867; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 200, 8)),
3 => std_logic_vector(to_unsigned( 37, 8)),
4 => std_logic_vector(to_unsigned( 214, 8)),
5 => std_logic_vector(to_unsigned( 40, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 196, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 24, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 12, 8)),
16 => std_logic_vector(to_unsigned( 246, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 199, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 867 then count <= 868; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 6, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 248, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 4, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 23, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 87, 8)),
11 => std_logic_vector(to_unsigned( 86, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 35, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 46, 8)),
18 => std_logic_vector(to_unsigned( 53, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 868 then count <= 869; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 196, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 32, 8)),
7 => std_logic_vector(to_unsigned( 102, 8)),
8 => std_logic_vector(to_unsigned( 36, 8)),
9 => std_logic_vector(to_unsigned( 184, 8)),
10 => std_logic_vector(to_unsigned( 56, 8)),
11 => std_logic_vector(to_unsigned( 92, 8)),
12 => std_logic_vector(to_unsigned( 201, 8)),
13 => std_logic_vector(to_unsigned( 155, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 29, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 869 then count <= 870; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 228, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 90, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 204, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 170, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 37, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 870 then count <= 871; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 189, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 253, 8)),
8 => std_logic_vector(to_unsigned( 239, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 178, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 172, 8)),
13 => std_logic_vector(to_unsigned( 94, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 45, 8)),
16 => std_logic_vector(to_unsigned( 191, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 871 then count <= 872; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 37, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 240, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 195, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 189, 8)),
9 => std_logic_vector(to_unsigned( 96, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 167, 8)),
12 => std_logic_vector(to_unsigned( 252, 8)),
13 => std_logic_vector(to_unsigned( 4, 8)),
14 => std_logic_vector(to_unsigned( 236, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 201, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 872 then count <= 873; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 21, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 18, 8)),
6 => std_logic_vector(to_unsigned( 184, 8)),
7 => std_logic_vector(to_unsigned( 10, 8)),
8 => std_logic_vector(to_unsigned( 29, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 71, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110010
elsif count = 873 then count <= 874; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 45, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 30, 8)),
4 => std_logic_vector(to_unsigned( 212, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 37, 8)),
7 => std_logic_vector(to_unsigned( 135, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 27, 8)),
12 => std_logic_vector(to_unsigned( 88, 8)),
13 => std_logic_vector(to_unsigned( 240, 8)),
14 => std_logic_vector(to_unsigned( 13, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 252, 8)),
17 => std_logic_vector(to_unsigned( 81, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 874 then count <= 875; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 50, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 36, 8)),
10 => std_logic_vector(to_unsigned( 18, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 18, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 50, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 875 then count <= 876; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 67, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 118, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 210, 8)),
8 => std_logic_vector(to_unsigned( 35, 8)),
9 => std_logic_vector(to_unsigned( 77, 8)),
10 => std_logic_vector(to_unsigned( 107, 8)),
11 => std_logic_vector(to_unsigned( 176, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 173, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 876 then count <= 877; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 39, 8)),
7 => std_logic_vector(to_unsigned( 195, 8)),
8 => std_logic_vector(to_unsigned( 91, 8)),
9 => std_logic_vector(to_unsigned( 226, 8)),
10 => std_logic_vector(to_unsigned( 4, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 230, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 231, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 205, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 877 then count <= 878; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 68, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 233, 8)),
5 => std_logic_vector(to_unsigned( 252, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 164, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 145, 8)),
10 => std_logic_vector(to_unsigned( 59, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 51, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 47, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011000
elsif count = 878 then count <= 879; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 25, 8)),
2 => std_logic_vector(to_unsigned( 84, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 241, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 8, 8)),
13 => std_logic_vector(to_unsigned( 15, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 49, 8)),
16 => std_logic_vector(to_unsigned( 132, 8)),
17 => std_logic_vector(to_unsigned( 53, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 879 then count <= 880; RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 118, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 155, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 42, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 17, 8)),
13 => std_logic_vector(to_unsigned( 170, 8)),
14 => std_logic_vector(to_unsigned( 181, 8)),
15 => std_logic_vector(to_unsigned( 172, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 880 then count <= 881; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 240, 8)),
4 => std_logic_vector(to_unsigned( 228, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 185, 8)),
7 => std_logic_vector(to_unsigned( 210, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 165, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 226, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 881 then count <= 882; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 86, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 230, 8)),
8 => std_logic_vector(to_unsigned( 3, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 73, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 80, 8)),
17 => std_logic_vector(to_unsigned( 54, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 882 then count <= 883; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 254, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 239, 8)),
4 => std_logic_vector(to_unsigned( 184, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 169, 8)),
9 => std_logic_vector(to_unsigned( 126, 8)),
10 => std_logic_vector(to_unsigned( 214, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 883 then count <= 884; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 62, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 27, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 74, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 119, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 88, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 126, 8)),
15 => std_logic_vector(to_unsigned( 251, 8)),
16 => std_logic_vector(to_unsigned( 249, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 884 then count <= 885; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 188, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 45, 8)),
5 => std_logic_vector(to_unsigned( 133, 8)),
6 => std_logic_vector(to_unsigned( 4, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 250, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 66, 8)),
12 => std_logic_vector(to_unsigned( 196, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 179, 8)),
15 => std_logic_vector(to_unsigned( 18, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 885 then count <= 886; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 45, 8)),
4 => std_logic_vector(to_unsigned( 2, 8)),
5 => std_logic_vector(to_unsigned( 226, 8)),
6 => std_logic_vector(to_unsigned( 60, 8)),
7 => std_logic_vector(to_unsigned( 218, 8)),
8 => std_logic_vector(to_unsigned( 52, 8)),
9 => std_logic_vector(to_unsigned( 66, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 204, 8)),
12 => std_logic_vector(to_unsigned( 44, 8)),
13 => std_logic_vector(to_unsigned( 220, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 56, 8)),
17 => std_logic_vector(to_unsigned( 207, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 886 then count <= 887; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 178, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 27, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 47, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 10, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 194, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 43, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 887 then count <= 888; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 116, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 159, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 23, 8)),
6 => std_logic_vector(to_unsigned( 193, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 74, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 14, 8)),
14 => std_logic_vector(to_unsigned( 239, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 888 then count <= 889; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 179, 8)),
6 => std_logic_vector(to_unsigned( 3, 8)),
7 => std_logic_vector(to_unsigned( 78, 8)),
8 => std_logic_vector(to_unsigned( 4, 8)),
9 => std_logic_vector(to_unsigned( 214, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 65, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 105, 8)),
15 => std_logic_vector(to_unsigned( 246, 8)),
16 => std_logic_vector(to_unsigned( 230, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 889 then count <= 890; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 183, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 176, 8)),
8 => std_logic_vector(to_unsigned( 56, 8)),
9 => std_logic_vector(to_unsigned( 12, 8)),
10 => std_logic_vector(to_unsigned( 175, 8)),
11 => std_logic_vector(to_unsigned( 48, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 155, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 890 then count <= 891; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 22, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 217, 8)),
5 => std_logic_vector(to_unsigned( 61, 8)),
6 => std_logic_vector(to_unsigned( 195, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 85, 8)),
12 => std_logic_vector(to_unsigned( 227, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 209, 8)),
15 => std_logic_vector(to_unsigned( 215, 8)),
16 => std_logic_vector(to_unsigned( 222, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 199, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 891 then count <= 892; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 145, 8)),
3 => std_logic_vector(to_unsigned( 50, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 52, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 238, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 22, 8)),
10 => std_logic_vector(to_unsigned( 229, 8)),
11 => std_logic_vector(to_unsigned( 236, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 78, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 892 then count <= 893; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 17, 8)),
5 => std_logic_vector(to_unsigned( 50, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 35, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 186, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 68, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 106, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 893 then count <= 894; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 129, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 246, 8)),
10 => std_logic_vector(to_unsigned( 112, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 135, 8)),
14 => std_logic_vector(to_unsigned( 135, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 894 then count <= 895; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 208, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 112, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 190, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 132, 8)),
12 => std_logic_vector(to_unsigned( 52, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 895 then count <= 896; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 204, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 18, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 48, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 28, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 33, 8)),
12 => std_logic_vector(to_unsigned( 59, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 45, 8)),
17 => std_logic_vector(to_unsigned( 53, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 896 then count <= 897; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 204, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 16, 8)),
5 => std_logic_vector(to_unsigned( 209, 8)),
6 => std_logic_vector(to_unsigned( 184, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 167, 8)),
12 => std_logic_vector(to_unsigned( 216, 8)),
13 => std_logic_vector(to_unsigned( 9, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 187, 8)),
16 => std_logic_vector(to_unsigned( 182, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 897 then count <= 898; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 246, 8)),
6 => std_logic_vector(to_unsigned( 67, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 92, 8)),
9 => std_logic_vector(to_unsigned( 213, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 164, 8)),
16 => std_logic_vector(to_unsigned( 225, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 898 then count <= 899; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 59, 8)),
4 => std_logic_vector(to_unsigned( 43, 8)),
5 => std_logic_vector(to_unsigned( 109, 8)),
6 => std_logic_vector(to_unsigned( 89, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 38, 8)),
10 => std_logic_vector(to_unsigned( 162, 8)),
11 => std_logic_vector(to_unsigned( 132, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 899 then count <= 900; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 8, 8)),
2 => std_logic_vector(to_unsigned( 61, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 26, 8)),
6 => std_logic_vector(to_unsigned( 252, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 247, 8)),
9 => std_logic_vector(to_unsigned( 99, 8)),
10 => std_logic_vector(to_unsigned( 237, 8)),
11 => std_logic_vector(to_unsigned( 112, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 136, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 105, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 900 then count <= 901; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 55, 8)),
2 => std_logic_vector(to_unsigned( 190, 8)),
3 => std_logic_vector(to_unsigned( 186, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 232, 8)),
7 => std_logic_vector(to_unsigned( 52, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 211, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 211, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 901 then count <= 902; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 249, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 92, 8)),
12 => std_logic_vector(to_unsigned( 160, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 0, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 902 then count <= 903; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 28, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 50, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 7, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 161, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 64, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 903 then count <= 904; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 3, 8)),
2 => std_logic_vector(to_unsigned( 207, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 47, 8)),
6 => std_logic_vector(to_unsigned( 230, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 83, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 78, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 904 then count <= 905; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 40, 8)),
4 => std_logic_vector(to_unsigned( 213, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 175, 8)),
7 => std_logic_vector(to_unsigned( 53, 8)),
8 => std_logic_vector(to_unsigned( 186, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 154, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 45, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 905 then count <= 906; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 218, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 193, 8)),
7 => std_logic_vector(to_unsigned( 255, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 46, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 250, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 198, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 80, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 906 then count <= 907; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 23, 8)),
2 => std_logic_vector(to_unsigned( 82, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 178, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 64, 8)),
8 => std_logic_vector(to_unsigned( 23, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 197, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 21, 8)),
15 => std_logic_vector(to_unsigned( 170, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 907 then count <= 908; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 217, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 84, 8)),
4 => std_logic_vector(to_unsigned( 241, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 233, 8)),
7 => std_logic_vector(to_unsigned( 85, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 76, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 34, 8)),
14 => std_logic_vector(to_unsigned( 182, 8)),
15 => std_logic_vector(to_unsigned( 32, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 908 then count <= 909; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 241, 8)),
3 => std_logic_vector(to_unsigned( 6, 8)),
4 => std_logic_vector(to_unsigned( 199, 8)),
5 => std_logic_vector(to_unsigned( 115, 8)),
6 => std_logic_vector(to_unsigned( 202, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 12, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 173, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 31, 8)),
14 => std_logic_vector(to_unsigned( 30, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00100111
elsif count = 909 then count <= 910; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 10, 8)),
4 => std_logic_vector(to_unsigned( 220, 8)),
5 => std_logic_vector(to_unsigned( 180, 8)),
6 => std_logic_vector(to_unsigned( 216, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 180, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 910 then count <= 911; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 136, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 205, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 71, 8)),
11 => std_logic_vector(to_unsigned( 214, 8)),
12 => std_logic_vector(to_unsigned( 244, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 28, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 911 then count <= 912; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 225, 8)),
3 => std_logic_vector(to_unsigned( 214, 8)),
4 => std_logic_vector(to_unsigned( 208, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 78, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 21, 8)),
11 => std_logic_vector(to_unsigned( 198, 8)),
12 => std_logic_vector(to_unsigned( 172, 8)),
13 => std_logic_vector(to_unsigned( 220, 8)),
14 => std_logic_vector(to_unsigned( 194, 8)),
15 => std_logic_vector(to_unsigned( 31, 8)),
16 => std_logic_vector(to_unsigned( 205, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 198, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 912 then count <= 913; RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 17, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 181, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 255, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 24, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 245, 8)),
12 => std_logic_vector(to_unsigned( 4, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 39, 8)),
17 => std_logic_vector(to_unsigned( 208, 8)),
18 => std_logic_vector(to_unsigned( 37, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 913 then count <= 914; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 60, 8)),
2 => std_logic_vector(to_unsigned( 202, 8)),
3 => std_logic_vector(to_unsigned( 182, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 251, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 167, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 46, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 177, 8)),
15 => std_logic_vector(to_unsigned( 228, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 53, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 914 then count <= 915; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 5, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 23, 8)),
5 => std_logic_vector(to_unsigned( 32, 8)),
6 => std_logic_vector(to_unsigned( 34, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 9, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 107, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 240, 8)),
14 => std_logic_vector(to_unsigned( 250, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 145, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 58, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 915 then count <= 916; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 25, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 195, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 151, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 244, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 916 then count <= 917; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 193, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 235, 8)),
6 => std_logic_vector(to_unsigned( 134, 8)),
7 => std_logic_vector(to_unsigned( 213, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 202, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 227, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 213, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 205, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 917 then count <= 918; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 220, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 246, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 112, 8)),
6 => std_logic_vector(to_unsigned( 1, 8)),
7 => std_logic_vector(to_unsigned( 237, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 179, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 243, 8)),
14 => std_logic_vector(to_unsigned( 116, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 156, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 918 then count <= 919; RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 220, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 100, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 241, 8)),
14 => std_logic_vector(to_unsigned( 231, 8)),
15 => std_logic_vector(to_unsigned( 226, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 919 then count <= 920; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 189, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 26, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 193, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110110
elsif count = 920 then count <= 921; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 51, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 29, 8)),
7 => std_logic_vector(to_unsigned( 3, 8)),
8 => std_logic_vector(to_unsigned( 153, 8)),
9 => std_logic_vector(to_unsigned( 36, 8)),
10 => std_logic_vector(to_unsigned( 2, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 59, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 921 then count <= 922; RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 139, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 34, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 229, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 56, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 234, 8)),
15 => std_logic_vector(to_unsigned( 152, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 922 then count <= 923; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 22, 8)),
3 => std_logic_vector(to_unsigned( 108, 8)),
4 => std_logic_vector(to_unsigned( 80, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 44, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 251, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 45, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 63, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 923 then count <= 924; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 62, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 90, 8)),
6 => std_logic_vector(to_unsigned( 159, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 28, 8)),
10 => std_logic_vector(to_unsigned( 178, 8)),
11 => std_logic_vector(to_unsigned( 216, 8)),
12 => std_logic_vector(to_unsigned( 180, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 88, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 924 then count <= 925; RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 54, 8)),
2 => std_logic_vector(to_unsigned( 253, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 203, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 237, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 227, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 188, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 144, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101100
elsif count = 925 then count <= 926; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 195, 8)),
2 => std_logic_vector(to_unsigned( 207, 8)),
3 => std_logic_vector(to_unsigned( 18, 8)),
4 => std_logic_vector(to_unsigned( 66, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 137, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 926 then count <= 927; RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 210, 8)),
3 => std_logic_vector(to_unsigned( 234, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 42, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 80, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110101
elsif count = 927 then count <= 928; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 208, 8)),
2 => std_logic_vector(to_unsigned( 112, 8)),
3 => std_logic_vector(to_unsigned( 23, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 189, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 199, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 77, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 928 then count <= 929; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 248, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 170, 8)),
6 => std_logic_vector(to_unsigned( 241, 8)),
7 => std_logic_vector(to_unsigned( 223, 8)),
8 => std_logic_vector(to_unsigned( 188, 8)),
9 => std_logic_vector(to_unsigned( 230, 8)),
10 => std_logic_vector(to_unsigned( 94, 8)),
11 => std_logic_vector(to_unsigned( 215, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 136, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 222, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 929 then count <= 930; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 165, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 108, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 32, 8)),
16 => std_logic_vector(to_unsigned( 98, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 930 then count <= 931; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 71, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 226, 8)),
5 => std_logic_vector(to_unsigned( 133, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 161, 8)),
8 => std_logic_vector(to_unsigned( 166, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 153, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 23, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 198, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 931 then count <= 932; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 82, 8)),
8 => std_logic_vector(to_unsigned( 245, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 19, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 51, 8)),
14 => std_logic_vector(to_unsigned( 214, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 245, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 210, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 932 then count <= 933; RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 50, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 48, 8)),
9 => std_logic_vector(to_unsigned( 224, 8)),
10 => std_logic_vector(to_unsigned( 44, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 188, 8)),
13 => std_logic_vector(to_unsigned( 250, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 90, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00100111
elsif count = 933 then count <= 934; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 241, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 248, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 183, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 116, 8)),
11 => std_logic_vector(to_unsigned( 172, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 20, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 213, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 934 then count <= 935; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 66, 8)),
2 => std_logic_vector(to_unsigned( 51, 8)),
3 => std_logic_vector(to_unsigned( 86, 8)),
4 => std_logic_vector(to_unsigned( 95, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 58, 8)),
9 => std_logic_vector(to_unsigned( 99, 8)),
10 => std_logic_vector(to_unsigned( 242, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 35, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 35, 8)),
15 => std_logic_vector(to_unsigned( 239, 8)),
16 => std_logic_vector(to_unsigned( 126, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 63, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 935 then count <= 936; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 31, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 45, 8)),
7 => std_logic_vector(to_unsigned( 214, 8)),
8 => std_logic_vector(to_unsigned( 100, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 13, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 936 then count <= 937; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 251, 8)),
2 => std_logic_vector(to_unsigned( 179, 8)),
3 => std_logic_vector(to_unsigned( 218, 8)),
4 => std_logic_vector(to_unsigned( 140, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 146, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 34, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 937 then count <= 938; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 195, 8)),
4 => std_logic_vector(to_unsigned( 91, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 210, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 25, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 249, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 938 then count <= 939; RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 120, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 170, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 156, 8)),
12 => std_logic_vector(to_unsigned( 116, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 139, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 939 then count <= 940; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 219, 8)),
4 => std_logic_vector(to_unsigned( 234, 8)),
5 => std_logic_vector(to_unsigned( 15, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 245, 8)),
9 => std_logic_vector(to_unsigned( 198, 8)),
10 => std_logic_vector(to_unsigned( 22, 8)),
11 => std_logic_vector(to_unsigned( 48, 8)),
12 => std_logic_vector(to_unsigned( 213, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 222, 8)),
15 => std_logic_vector(to_unsigned( 61, 8)),
16 => std_logic_vector(to_unsigned( 226, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 940 then count <= 941; RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 62, 8)),
4 => std_logic_vector(to_unsigned( 32, 8)),
5 => std_logic_vector(to_unsigned( 205, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 57, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 172, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 941 then count <= 942; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 48, 8)),
3 => std_logic_vector(to_unsigned( 190, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 218, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 46, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 9, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 942 then count <= 943; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 157, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 205, 8)),
5 => std_logic_vector(to_unsigned( 232, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 206, 8)),
9 => std_logic_vector(to_unsigned( 156, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 0, 8)),
12 => std_logic_vector(to_unsigned( 57, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 73, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 943 then count <= 944; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 219, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 192, 8)),
6 => std_logic_vector(to_unsigned( 243, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 111, 8)),
10 => std_logic_vector(to_unsigned( 207, 8)),
11 => std_logic_vector(to_unsigned( 112, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 944 then count <= 945; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 55, 8)),
3 => std_logic_vector(to_unsigned( 194, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 177, 8)),
10 => std_logic_vector(to_unsigned( 51, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 85, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 242, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 189, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 945 then count <= 946; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 21, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 58, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 69, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 255, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 47, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101100
elsif count = 946 then count <= 947; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 232, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 47, 8)),
6 => std_logic_vector(to_unsigned( 83, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 6, 8)),
9 => std_logic_vector(to_unsigned( 72, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 76, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 947 then count <= 948; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 55, 8)),
2 => std_logic_vector(to_unsigned( 193, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 181, 8)),
5 => std_logic_vector(to_unsigned( 110, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 251, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 177, 8)),
13 => std_logic_vector(to_unsigned( 87, 8)),
14 => std_logic_vector(to_unsigned( 26, 8)),
15 => std_logic_vector(to_unsigned( 78, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 190, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 948 then count <= 949; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 17, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 146, 8)),
6 => std_logic_vector(to_unsigned( 54, 8)),
7 => std_logic_vector(to_unsigned( 188, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 35, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 173, 8)),
13 => std_logic_vector(to_unsigned( 226, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 949 then count <= 950; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 143, 8)),
3 => std_logic_vector(to_unsigned( 4, 8)),
4 => std_logic_vector(to_unsigned( 77, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 25, 8)),
10 => std_logic_vector(to_unsigned( 8, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 212, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 141, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 950 then count <= 951; RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 232, 8)),
3 => std_logic_vector(to_unsigned( 178, 8)),
4 => std_logic_vector(to_unsigned( 250, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 186, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 226, 8)),
13 => std_logic_vector(to_unsigned( 170, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 247, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 221, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 951 then count <= 952; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 245, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 241, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 112, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 229, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 197, 8)),
14 => std_logic_vector(to_unsigned( 140, 8)),
15 => std_logic_vector(to_unsigned( 9, 8)),
16 => std_logic_vector(to_unsigned( 51, 8)),
17 => std_logic_vector(to_unsigned( 223, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 952 then count <= 953; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 228, 8)),
2 => std_logic_vector(to_unsigned( 112, 8)),
3 => std_logic_vector(to_unsigned( 48, 8)),
4 => std_logic_vector(to_unsigned( 50, 8)),
5 => std_logic_vector(to_unsigned( 51, 8)),
6 => std_logic_vector(to_unsigned( 66, 8)),
7 => std_logic_vector(to_unsigned( 44, 8)),
8 => std_logic_vector(to_unsigned( 248, 8)),
9 => std_logic_vector(to_unsigned( 226, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 210, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 175, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 221, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 953 then count <= 954; RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 52, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 116, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 954 then count <= 955; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 31, 8)),
2 => std_logic_vector(to_unsigned( 227, 8)),
3 => std_logic_vector(to_unsigned( 28, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 86, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 85, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 78, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 69, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 105, 8)),
17 => std_logic_vector(to_unsigned( 118, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 955 then count <= 956; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 209, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 214, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 197, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 2, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 119, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 20, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 956 then count <= 957; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 187, 8)),
3 => std_logic_vector(to_unsigned( 12, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 230, 8)),
6 => std_logic_vector(to_unsigned( 17, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 36, 8)),
9 => std_logic_vector(to_unsigned( 33, 8)),
10 => std_logic_vector(to_unsigned( 142, 8)),
11 => std_logic_vector(to_unsigned( 6, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 39, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 63, 8)),
16 => std_logic_vector(to_unsigned( 210, 8)),
17 => std_logic_vector(to_unsigned( 55, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 957 then count <= 958; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 248, 8)),
2 => std_logic_vector(to_unsigned( 3, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 9, 8)),
5 => std_logic_vector(to_unsigned( 61, 8)),
6 => std_logic_vector(to_unsigned( 159, 8)),
7 => std_logic_vector(to_unsigned( 38, 8)),
8 => std_logic_vector(to_unsigned( 21, 8)),
9 => std_logic_vector(to_unsigned( 58, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 32, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100100
elsif count = 958 then count <= 959; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 87, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 233, 8)),
6 => std_logic_vector(to_unsigned( 62, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 149, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 36, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 241, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 190, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011010
elsif count = 959 then count <= 960; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 170, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 182, 8)),
7 => std_logic_vector(to_unsigned( 21, 8)),
8 => std_logic_vector(to_unsigned( 0, 8)),
9 => std_logic_vector(to_unsigned( 246, 8)),
10 => std_logic_vector(to_unsigned( 60, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 186, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 960 then count <= 961; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 205, 8)),
2 => std_logic_vector(to_unsigned( 142, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 109, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 189, 8)),
9 => std_logic_vector(to_unsigned( 215, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 37, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 57, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 197, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 961 then count <= 962; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 252, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 219, 8)),
4 => std_logic_vector(to_unsigned( 155, 8)),
5 => std_logic_vector(to_unsigned( 115, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 199, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 76, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 180, 8)),
13 => std_logic_vector(to_unsigned( 135, 8)),
14 => std_logic_vector(to_unsigned( 244, 8)),
15 => std_logic_vector(to_unsigned( 197, 8)),
16 => std_logic_vector(to_unsigned( 185, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100110
elsif count = 962 then count <= 963; RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 239, 8)),
2 => std_logic_vector(to_unsigned( 209, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 222, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 200, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 75, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 46, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 963 then count <= 964; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 199, 8)),
5 => std_logic_vector(to_unsigned( 229, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 183, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 218, 8)),
16 => std_logic_vector(to_unsigned( 162, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 964 then count <= 965; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 78, 8)),
2 => std_logic_vector(to_unsigned( 192, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 207, 8)),
7 => std_logic_vector(to_unsigned( 77, 8)),
8 => std_logic_vector(to_unsigned( 191, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 45, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 965 then count <= 966; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 65, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 133, 8)),
6 => std_logic_vector(to_unsigned( 231, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 227, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 31, 8)),
12 => std_logic_vector(to_unsigned( 35, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 214, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 210, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 966 then count <= 967; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 1, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 153, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 237, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 116, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 34, 8)),
11 => std_logic_vector(to_unsigned( 150, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 245, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 53, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 967 then count <= 968; RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 71, 8)),
3 => std_logic_vector(to_unsigned( 81, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 207, 8)),
7 => std_logic_vector(to_unsigned( 150, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 23, 8)),
10 => std_logic_vector(to_unsigned( 246, 8)),
11 => std_logic_vector(to_unsigned( 192, 8)),
12 => std_logic_vector(to_unsigned( 34, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 204, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 191, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 203, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 968 then count <= 969; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 156, 8)),
3 => std_logic_vector(to_unsigned( 200, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 31, 8)),
6 => std_logic_vector(to_unsigned( 251, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 15, 8)),
9 => std_logic_vector(to_unsigned( 76, 8)),
10 => std_logic_vector(to_unsigned( 252, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 969 then count <= 970; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 9, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 132, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 117, 8)),
11 => std_logic_vector(to_unsigned( 209, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 184, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 970 then count <= 971; RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 60, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 158, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 165, 8)),
11 => std_logic_vector(to_unsigned( 183, 8)),
12 => std_logic_vector(to_unsigned( 244, 8)),
13 => std_logic_vector(to_unsigned( 152, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 193, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 971 then count <= 972; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 221, 8)),
2 => std_logic_vector(to_unsigned( 222, 8)),
3 => std_logic_vector(to_unsigned( 112, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 60, 8)),
7 => std_logic_vector(to_unsigned( 237, 8)),
8 => std_logic_vector(to_unsigned( 206, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 13, 8)),
11 => std_logic_vector(to_unsigned( 172, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 236, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 5, 8)),
17 => std_logic_vector(to_unsigned( 204, 8)),
18 => std_logic_vector(to_unsigned( 206, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 972 then count <= 973; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 168, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 101, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 38, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 242, 8)),
8 => std_logic_vector(to_unsigned( 61, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 9, 8)),
13 => std_logic_vector(to_unsigned( 22, 8)),
14 => std_logic_vector(to_unsigned( 215, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 59, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 973 then count <= 974; RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 155, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 59, 8)),
6 => std_logic_vector(to_unsigned( 89, 8)),
7 => std_logic_vector(to_unsigned( 254, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 184, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 229, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 974 then count <= 975; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 19, 8)),
2 => std_logic_vector(to_unsigned( 42, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 161, 8)),
6 => std_logic_vector(to_unsigned( 231, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 94, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 243, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 975 then count <= 976; RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 55, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 70, 8)),
11 => std_logic_vector(to_unsigned( 95, 8)),
12 => std_logic_vector(to_unsigned( 201, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 79, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 976 then count <= 977; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 209, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 231, 8)),
5 => std_logic_vector(to_unsigned( 122, 8)),
6 => std_logic_vector(to_unsigned( 66, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 12, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 193, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101100
elsif count = 977 then count <= 978; RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 24, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 180, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 179, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 978 then count <= 979; RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 127, 8)),
4 => std_logic_vector(to_unsigned( 73, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 67, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 200, 8)),
10 => std_logic_vector(to_unsigned( 16, 8)),
11 => std_logic_vector(to_unsigned( 243, 8)),
12 => std_logic_vector(to_unsigned( 253, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 979 then count <= 980; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 207, 8)),
5 => std_logic_vector(to_unsigned( 101, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 21, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 76, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 980 then count <= 981; RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 170, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 49, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 30, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 247, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 231, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 12, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 981 then count <= 982; RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 195, 8)),
4 => std_logic_vector(to_unsigned( 233, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 89, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 184, 8)),
12 => std_logic_vector(to_unsigned( 71, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 63, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 982 then count <= 983; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 187, 8)),
3 => std_logic_vector(to_unsigned( 100, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 207, 8)),
7 => std_logic_vector(to_unsigned( 211, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 99, 8)),
10 => std_logic_vector(to_unsigned( 221, 8)),
11 => std_logic_vector(to_unsigned( 224, 8)),
12 => std_logic_vector(to_unsigned( 34, 8)),
13 => std_logic_vector(to_unsigned( 87, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 38, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 190, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 983 then count <= 984; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 221, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 233, 8)),
5 => std_logic_vector(to_unsigned( 77, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 249, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 122, 8)),
11 => std_logic_vector(to_unsigned( 226, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 235, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 984 then count <= 985; RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 191, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 78, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 112, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 48, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 42, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 985 then count <= 986; RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 196, 8)),
2 => std_logic_vector(to_unsigned( 91, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 19, 8)),
12 => std_logic_vector(to_unsigned( 84, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 46, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 986 then count <= 987; RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 163, 8)),
2 => std_logic_vector(to_unsigned( 36, 8)),
3 => std_logic_vector(to_unsigned( 56, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 111, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 26, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 91, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110110
elsif count = 987 then count <= 988; RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 192, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 29, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 988 then count <= 989; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 177, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 204, 8)),
4 => std_logic_vector(to_unsigned( 95, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 41, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 230, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 225, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 989 then count <= 990; RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 55, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 59, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 147, 8)),
8 => std_logic_vector(to_unsigned( 151, 8)),
9 => std_logic_vector(to_unsigned( 42, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 205, 8)),
12 => std_logic_vector(to_unsigned( 2, 8)),
13 => std_logic_vector(to_unsigned( 178, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 57, 8)),
16 => std_logic_vector(to_unsigned( 83, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 990 then count <= 991; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 208, 8)),
2 => std_logic_vector(to_unsigned( 219, 8)),
3 => std_logic_vector(to_unsigned( 91, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 4, 8)),
12 => std_logic_vector(to_unsigned( 75, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 237, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 185, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 991 then count <= 992; RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 22, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 33, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 37, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 0, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 47, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 28, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 249, 8)),
15 => std_logic_vector(to_unsigned( 25, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 76, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 992 then count <= 993; RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 92, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 186, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 241, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 993 then count <= 994; RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 176, 8)),
8 => std_logic_vector(to_unsigned( 130, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 13, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 994 then count <= 995; RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 22, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 55, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 198, 8)),
7 => std_logic_vector(to_unsigned( 148, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 185, 8)),
13 => std_logic_vector(to_unsigned( 254, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 995 then count <= 996; RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 3, 8)),
2 => std_logic_vector(to_unsigned( 4, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 4, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 134, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 36, 8)),
12 => std_logic_vector(to_unsigned( 110, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 58, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 996 then count <= 997; RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 228, 8)),
2 => std_logic_vector(to_unsigned( 41, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 123, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 166, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 106, 8)),
9 => std_logic_vector(to_unsigned( 239, 8)),
10 => std_logic_vector(to_unsigned( 8, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 45, 8)),
15 => std_logic_vector(to_unsigned( 33, 8)),
16 => std_logic_vector(to_unsigned( 182, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101110
elsif count = 997 then count <= 998; RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 60, 8)),
2 => std_logic_vector(to_unsigned( 72, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 243, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 32, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 998 then count <= 999; RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 148, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 14, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 86, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 8, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 207, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 999 then count <= 1000; RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 94, 8)),
2 => std_logic_vector(to_unsigned( 218, 8)),
3 => std_logic_vector(to_unsigned( 1, 8)),
4 => std_logic_vector(to_unsigned( 18, 8)),
5 => std_logic_vector(to_unsigned( 23, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 100, 8)),
9 => std_logic_vector(to_unsigned( 96, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 34, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 250, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001101
end if; end if;
                end process;
                test : process is
                begin wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101110" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001101" report "TEST FAILED" severity failure;assert false report "1000 TESTS PASSED" severity failure;
    end process test;
                end projecttb;