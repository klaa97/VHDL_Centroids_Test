library ieee;
                use ieee.std_logic_1164.all;
                use ieee.numeric_std.all;
                use ieee.std_logic_unsigned.all;
                entity multiple_test is
                end multiple_test;
                architecture projecttb of multiple_test is
                constant c_CLOCK_PERIOD		: time := 100 ns;
                signal   tb_done		: std_logic;
                signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
                signal   tb_rst	                : std_logic := '0';
                signal   tb_start		: std_logic := '0';
                signal   tb_clk		        : std_logic := '0';
                signal   mem_o_data,mem_i_data	: std_logic_vector (7 downto 0);
                signal   enable_wire  		: std_logic;
                signal   mem_we		        : std_logic;
                type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
                signal RAM: ram_type := (0 => "11101110",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 232, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 224, 8)),
7 => std_logic_vector(to_unsigned( 213, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 51, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 200, 8)),
 others => (others => '0'));
signal count : integer := 0;
-- MASK_OUT: 	 10101110
 component project_reti_logiche is
                port (
                    i_clk         : in  std_logic;
                    i_start       : in  std_logic;
                    i_rst         : in  std_logic;
                    i_data        : in  std_logic_vector(7 downto 0);
                    o_address     : out std_logic_vector(15 downto 0);
                    o_done        : out std_logic;
                    o_en          : out std_logic;
                    o_we          : out std_logic;
                    o_data        : out std_logic_vector (7 downto 0)
                    );
                end component project_reti_logiche;
                begin
                UUT: project_reti_logiche
                port map (
                        i_clk      	=> tb_clk,
                        i_start       => tb_start,
                        i_rst      	=> tb_rst,
                        i_data    	=> mem_o_data,
                        o_address  	=> mem_address,
                        o_done      	=> tb_done,
                        o_en   	=> enable_wire,
                        o_we 		=> mem_we,
                        o_data    	=> mem_i_data
                        );
                p_CLK_GEN : process is
                begin
                    wait for c_CLOCK_PERIOD/2;
                    tb_clk <= not tb_clk;
                end process p_CLK_GEN;
                MEM : process(tb_clk)
                begin
                    if tb_clk'event and tb_clk = '1' then
                        if enable_wire = '1' then
                            if mem_we = '1' then
                                RAM(conv_integer(mem_address))  <= mem_i_data;
                                mem_o_data                      <= mem_i_data after 2 ns;
                            else
                                mem_o_data <= RAM(conv_integer(mem_address)) after 2 ns;
                            end if;
                        end if;
                    else if count = 1 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 216, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 45, 8)),
5 => std_logic_vector(to_unsigned( 181, 8)),
6 => std_logic_vector(to_unsigned( 62, 8)),
7 => std_logic_vector(to_unsigned( 173, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 208, 8)),
10 => std_logic_vector(to_unsigned( 119, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 58, 8)),
13 => std_logic_vector(to_unsigned( 218, 8)),
14 => std_logic_vector(to_unsigned( 57, 8)),
15 => std_logic_vector(to_unsigned( 241, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 202, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 2 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 61, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 64, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 145, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 3 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 42, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 20, 8)),
5 => std_logic_vector(to_unsigned( 41, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 65, 8)),
9 => std_logic_vector(to_unsigned( 177, 8)),
10 => std_logic_vector(to_unsigned( 11, 8)),
11 => std_logic_vector(to_unsigned( 199, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 180, 8)),
15 => std_logic_vector(to_unsigned( 68, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 4 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 99, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 249, 8)),
4 => std_logic_vector(to_unsigned( 207, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 114, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 106, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 161, 8)),
12 => std_logic_vector(to_unsigned( 0, 8)),
13 => std_logic_vector(to_unsigned( 157, 8)),
14 => std_logic_vector(to_unsigned( 85, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 5 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 203, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 161, 8)),
8 => std_logic_vector(to_unsigned( 13, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 58, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 6 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 7, 8)),
4 => std_logic_vector(to_unsigned( 199, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 199, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 38, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 90, 8)),
15 => std_logic_vector(to_unsigned( 113, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 7 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 229, 8)),
3 => std_logic_vector(to_unsigned( 216, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 218, 8)),
6 => std_logic_vector(to_unsigned( 184, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 230, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 221, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 94, 8)),
14 => std_logic_vector(to_unsigned( 211, 8)),
15 => std_logic_vector(to_unsigned( 56, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 8 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 188, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 232, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 178, 8)),
7 => std_logic_vector(to_unsigned( 154, 8)),
8 => std_logic_vector(to_unsigned( 235, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 29, 8)),
13 => std_logic_vector(to_unsigned( 221, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 159, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 203, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 9 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 149, 8)),
4 => std_logic_vector(to_unsigned( 16, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 37, 8)),
8 => std_logic_vector(to_unsigned( 207, 8)),
9 => std_logic_vector(to_unsigned( 182, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 214, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 149, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110101
elsif count = 10 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 205, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 175, 8)),
7 => std_logic_vector(to_unsigned( 135, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 19, 8)),
11 => std_logic_vector(to_unsigned( 231, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 224, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 11 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 216, 8)),
5 => std_logic_vector(to_unsigned( 198, 8)),
6 => std_logic_vector(to_unsigned( 202, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 239, 8)),
11 => std_logic_vector(to_unsigned( 191, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 33, 8)),
14 => std_logic_vector(to_unsigned( 231, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 218, 8)),
18 => std_logic_vector(to_unsigned( 185, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 12 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 130, 8)),
3 => std_logic_vector(to_unsigned( 21, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 110, 8)),
6 => std_logic_vector(to_unsigned( 204, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 64, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 22, 8)),
13 => std_logic_vector(to_unsigned( 56, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 250, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 13 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 233, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 47, 8)),
5 => std_logic_vector(to_unsigned( 134, 8)),
6 => std_logic_vector(to_unsigned( 208, 8)),
7 => std_logic_vector(to_unsigned( 10, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 216, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 186, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 181, 8)),
18 => std_logic_vector(to_unsigned( 200, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 14 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 29, 8)),
3 => std_logic_vector(to_unsigned( 56, 8)),
4 => std_logic_vector(to_unsigned( 74, 8)),
5 => std_logic_vector(to_unsigned( 78, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 54, 8)),
8 => std_logic_vector(to_unsigned( 78, 8)),
9 => std_logic_vector(to_unsigned( 244, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 29, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 15 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 39, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 36, 8)),
6 => std_logic_vector(to_unsigned( 166, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 74, 8)),
10 => std_logic_vector(to_unsigned( 250, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 229, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 28, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 145, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 16 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 54, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 7, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 161, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 214, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 161, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 240, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 17 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 95, 8)),
2 => std_logic_vector(to_unsigned( 177, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 187, 8)),
5 => std_logic_vector(to_unsigned( 41, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 144, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 136, 8)),
12 => std_logic_vector(to_unsigned( 198, 8)),
13 => std_logic_vector(to_unsigned( 178, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 61, 8)),
16 => std_logic_vector(to_unsigned( 170, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 18 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 113, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 155, 8)),
16 => std_logic_vector(to_unsigned( 15, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 19 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 25, 8)),
4 => std_logic_vector(to_unsigned( 50, 8)),
5 => std_logic_vector(to_unsigned( 115, 8)),
6 => std_logic_vector(to_unsigned( 66, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 20 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 62, 8)),
2 => std_logic_vector(to_unsigned( 233, 8)),
3 => std_logic_vector(to_unsigned( 197, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 163, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 204, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 100, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 88, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 21 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 10, 8)),
4 => std_logic_vector(to_unsigned( 181, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 211, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 203, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 240, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 22 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 240, 8)),
4 => std_logic_vector(to_unsigned( 99, 8)),
5 => std_logic_vector(to_unsigned( 93, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 166, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 64, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 200, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010011
elsif count = 23 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 19, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 102, 8)),
8 => std_logic_vector(to_unsigned( 34, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 212, 8)),
11 => std_logic_vector(to_unsigned( 28, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010101
elsif count = 24 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 39, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 35, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 120, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 210, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 25 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 202, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 182, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 145, 8)),
10 => std_logic_vector(to_unsigned( 243, 8)),
11 => std_logic_vector(to_unsigned( 167, 8)),
12 => std_logic_vector(to_unsigned( 18, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 37, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 244, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 26 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 23, 8)),
3 => std_logic_vector(to_unsigned( 169, 8)),
4 => std_logic_vector(to_unsigned( 74, 8)),
5 => std_logic_vector(to_unsigned( 47, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 47, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 83, 8)),
16 => std_logic_vector(to_unsigned( 191, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 27 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 112, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 221, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 28, 8)),
14 => std_logic_vector(to_unsigned( 69, 8)),
15 => std_logic_vector(to_unsigned( 245, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110101
elsif count = 28 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 94, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 5, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 76, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 28, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 40, 8)),
17 => std_logic_vector(to_unsigned( 76, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 29 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 85, 8)),
6 => std_logic_vector(to_unsigned( 81, 8)),
7 => std_logic_vector(to_unsigned( 39, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 215, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 30 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 211, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 227, 8)),
8 => std_logic_vector(to_unsigned( 92, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 221, 8)),
12 => std_logic_vector(to_unsigned( 86, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 253, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 80, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 31 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 33, 8)),
2 => std_logic_vector(to_unsigned( 94, 8)),
3 => std_logic_vector(to_unsigned( 47, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 58, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 32 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 42, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 226, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 75, 8)),
11 => std_logic_vector(to_unsigned( 55, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 55, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 81, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 33 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 87, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 216, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 203, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 34 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 219, 8)),
5 => std_logic_vector(to_unsigned( 44, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 66, 8)),
8 => std_logic_vector(to_unsigned( 140, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 156, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 36, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 35 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 233, 8)),
3 => std_logic_vector(to_unsigned( 76, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 92, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 74, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 51, 8)),
17 => std_logic_vector(to_unsigned( 48, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 36 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 243, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 1, 8)),
5 => std_logic_vector(to_unsigned( 26, 8)),
6 => std_logic_vector(to_unsigned( 219, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 206, 8)),
11 => std_logic_vector(to_unsigned( 112, 8)),
12 => std_logic_vector(to_unsigned( 189, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 18, 8)),
15 => std_logic_vector(to_unsigned( 164, 8)),
16 => std_logic_vector(to_unsigned( 195, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 203, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 37 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 221, 8)),
2 => std_logic_vector(to_unsigned( 34, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 13, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 245, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 62, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 51, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 38 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 166, 8)),
5 => std_logic_vector(to_unsigned( 192, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 196, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 39 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 117, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 44, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 146, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 85, 8)),
12 => std_logic_vector(to_unsigned( 204, 8)),
13 => std_logic_vector(to_unsigned( 6, 8)),
14 => std_logic_vector(to_unsigned( 252, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010110
elsif count = 40 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 49, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 209, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 184, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 219, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 222, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 41 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 20, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 240, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 48, 8)),
8 => std_logic_vector(to_unsigned( 230, 8)),
9 => std_logic_vector(to_unsigned( 15, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 29, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 126, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 55, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 42 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 206, 8)),
3 => std_logic_vector(to_unsigned( 65, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 51, 8)),
9 => std_logic_vector(to_unsigned( 81, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 253, 8)),
12 => std_logic_vector(to_unsigned( 7, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 66, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 53, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 43 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 24, 8)),
3 => std_logic_vector(to_unsigned( 165, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 51, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 177, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 178, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 191, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 138, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 44 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 180, 8)),
2 => std_logic_vector(to_unsigned( 182, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 118, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 51, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 198, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 45 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 171, 8)),
3 => std_logic_vector(to_unsigned( 27, 8)),
4 => std_logic_vector(to_unsigned( 219, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 62, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 106, 8)),
9 => std_logic_vector(to_unsigned( 110, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 219, 8)),
14 => std_logic_vector(to_unsigned( 205, 8)),
15 => std_logic_vector(to_unsigned( 104, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 46 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 152, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 62, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 2, 8)),
11 => std_logic_vector(to_unsigned( 37, 8)),
12 => std_logic_vector(to_unsigned( 151, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 30, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 47 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 173, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 133, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 155, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 48 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 229, 8)),
2 => std_logic_vector(to_unsigned( 236, 8)),
3 => std_logic_vector(to_unsigned( 201, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 220, 8)),
6 => std_logic_vector(to_unsigned( 245, 8)),
7 => std_logic_vector(to_unsigned( 150, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 210, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 31, 8)),
14 => std_logic_vector(to_unsigned( 83, 8)),
15 => std_logic_vector(to_unsigned( 230, 8)),
16 => std_logic_vector(to_unsigned( 235, 8)),
17 => std_logic_vector(to_unsigned( 210, 8)),
18 => std_logic_vector(to_unsigned( 221, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 49 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 197, 8)),
3 => std_logic_vector(to_unsigned( 75, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 98, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 48, 8)),
13 => std_logic_vector(to_unsigned( 35, 8)),
14 => std_logic_vector(to_unsigned( 7, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 50 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 175, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 227, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 41, 8)),
12 => std_logic_vector(to_unsigned( 216, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 51 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 168, 8)),
2 => std_logic_vector(to_unsigned( 240, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 248, 8)),
5 => std_logic_vector(to_unsigned( 37, 8)),
6 => std_logic_vector(to_unsigned( 8, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 247, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 18, 8)),
15 => std_logic_vector(to_unsigned( 253, 8)),
16 => std_logic_vector(to_unsigned( 131, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 52 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 4, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 212, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 199, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 53 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 165, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 165, 8)),
4 => std_logic_vector(to_unsigned( 214, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 127, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 238, 8)),
10 => std_logic_vector(to_unsigned( 23, 8)),
11 => std_logic_vector(to_unsigned( 173, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 208, 8)),
14 => std_logic_vector(to_unsigned( 82, 8)),
15 => std_logic_vector(to_unsigned( 252, 8)),
16 => std_logic_vector(to_unsigned( 3, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 54 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 91, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 184, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 248, 8)),
10 => std_logic_vector(to_unsigned( 24, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 56, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 55 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 51, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 10, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 28, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 201, 8)),
9 => std_logic_vector(to_unsigned( 3, 8)),
10 => std_logic_vector(to_unsigned( 44, 8)),
11 => std_logic_vector(to_unsigned( 41, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 9, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 244, 8)),
17 => std_logic_vector(to_unsigned( 44, 8)),
18 => std_logic_vector(to_unsigned( 44, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 56 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 215, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 37, 8)),
7 => std_logic_vector(to_unsigned( 204, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 136, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 235, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 230, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 242, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 210, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 57 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 91, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 74, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 148, 8)),
8 => std_logic_vector(to_unsigned( 28, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 83, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 58 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 168, 8)),
2 => std_logic_vector(to_unsigned( 130, 8)),
3 => std_logic_vector(to_unsigned( 196, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 90, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 217, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 63, 8)),
13 => std_logic_vector(to_unsigned( 224, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 90, 8)),
16 => std_logic_vector(to_unsigned( 236, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 59 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 74, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 47, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 136, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 21, 8)),
14 => std_logic_vector(to_unsigned( 135, 8)),
15 => std_logic_vector(to_unsigned( 36, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 73, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 60 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 252, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 225, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 237, 8)),
14 => std_logic_vector(to_unsigned( 172, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 61 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 60, 8)),
3 => std_logic_vector(to_unsigned( 35, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 76, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 212, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 8, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 62 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 149, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 78, 8)),
6 => std_logic_vector(to_unsigned( 103, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 119, 8)),
10 => std_logic_vector(to_unsigned( 216, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 11, 8)),
15 => std_logic_vector(to_unsigned( 132, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 63 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 220, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 245, 8)),
4 => std_logic_vector(to_unsigned( 235, 8)),
5 => std_logic_vector(to_unsigned( 240, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 190, 8)),
10 => std_logic_vector(to_unsigned( 9, 8)),
11 => std_logic_vector(to_unsigned( 65, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 204, 8)),
14 => std_logic_vector(to_unsigned( 50, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 78, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 64 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 41, 8)),
8 => std_logic_vector(to_unsigned( 204, 8)),
9 => std_logic_vector(to_unsigned( 76, 8)),
10 => std_logic_vector(to_unsigned( 255, 8)),
11 => std_logic_vector(to_unsigned( 210, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 211, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 65 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 214, 8)),
5 => std_logic_vector(to_unsigned( 124, 8)),
6 => std_logic_vector(to_unsigned( 227, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 214, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 232, 8)),
11 => std_logic_vector(to_unsigned( 203, 8)),
12 => std_logic_vector(to_unsigned( 12, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 177, 8)),
15 => std_logic_vector(to_unsigned( 123, 8)),
16 => std_logic_vector(to_unsigned( 190, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 209, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 66 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 76, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 191, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 215, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 223, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110010
elsif count = 67 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 247, 8)),
4 => std_logic_vector(to_unsigned( 235, 8)),
5 => std_logic_vector(to_unsigned( 170, 8)),
6 => std_logic_vector(to_unsigned( 31, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 79, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 251, 8)),
15 => std_logic_vector(to_unsigned( 132, 8)),
16 => std_logic_vector(to_unsigned( 178, 8)),
17 => std_logic_vector(to_unsigned( 44, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 68 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 61, 8)),
2 => std_logic_vector(to_unsigned( 57, 8)),
3 => std_logic_vector(to_unsigned( 28, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 32, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 41, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 9, 8)),
14 => std_logic_vector(to_unsigned( 249, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 44, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 69 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 212, 8)),
5 => std_logic_vector(to_unsigned( 233, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 119, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 132, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 70 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 230, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 88, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 56, 8)),
8 => std_logic_vector(to_unsigned( 61, 8)),
9 => std_logic_vector(to_unsigned( 170, 8)),
10 => std_logic_vector(to_unsigned( 230, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 16, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 60, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 71 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 148, 8)),
7 => std_logic_vector(to_unsigned( 9, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 41, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 161, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 15, 8)),
14 => std_logic_vector(to_unsigned( 83, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 72 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 153, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 86, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 60, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 68, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 126, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 73 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 170, 8)),
2 => std_logic_vector(to_unsigned( 94, 8)),
3 => std_logic_vector(to_unsigned( 255, 8)),
4 => std_logic_vector(to_unsigned( 99, 8)),
5 => std_logic_vector(to_unsigned( 42, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 230, 8)),
10 => std_logic_vector(to_unsigned( 116, 8)),
11 => std_logic_vector(to_unsigned( 31, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 212, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 74 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 44, 8)),
2 => std_logic_vector(to_unsigned( 131, 8)),
3 => std_logic_vector(to_unsigned( 171, 8)),
4 => std_logic_vector(to_unsigned( 243, 8)),
5 => std_logic_vector(to_unsigned( 36, 8)),
6 => std_logic_vector(to_unsigned( 239, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 209, 8)),
9 => std_logic_vector(to_unsigned( 5, 8)),
10 => std_logic_vector(to_unsigned( 212, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 216, 8)),
14 => std_logic_vector(to_unsigned( 138, 8)),
15 => std_logic_vector(to_unsigned( 194, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 75 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 230, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 228, 8)),
8 => std_logic_vector(to_unsigned( 207, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 129, 8)),
12 => std_logic_vector(to_unsigned( 43, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 78, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 76 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 158, 8)),
2 => std_logic_vector(to_unsigned( 23, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 220, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 73, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 76, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001010
elsif count = 77 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 53, 8)),
3 => std_logic_vector(to_unsigned( 7, 8)),
4 => std_logic_vector(to_unsigned( 249, 8)),
5 => std_logic_vector(to_unsigned( 190, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 103, 8)),
8 => std_logic_vector(to_unsigned( 75, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 205, 8)),
12 => std_logic_vector(to_unsigned( 85, 8)),
13 => std_logic_vector(to_unsigned( 181, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 167, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 78 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 254, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 43, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 32, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 30, 8)),
12 => std_logic_vector(to_unsigned( 90, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 72, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 79 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 211, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 35, 8)),
8 => std_logic_vector(to_unsigned( 59, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 80 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 89, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 230, 8)),
14 => std_logic_vector(to_unsigned( 30, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 81 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 58, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 48, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 25, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 66, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 48, 8)),
12 => std_logic_vector(to_unsigned( 222, 8)),
13 => std_logic_vector(to_unsigned( 173, 8)),
14 => std_logic_vector(to_unsigned( 31, 8)),
15 => std_logic_vector(to_unsigned( 80, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 46, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 82 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 210, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 9, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 220, 8)),
8 => std_logic_vector(to_unsigned( 24, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 10, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 187, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 177, 8)),
16 => std_logic_vector(to_unsigned( 132, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 83 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 166, 8)),
2 => std_logic_vector(to_unsigned( 228, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 8, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 163, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 99, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 84 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 55, 8)),
3 => std_logic_vector(to_unsigned( 113, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 222, 8)),
8 => std_logic_vector(to_unsigned( 106, 8)),
9 => std_logic_vector(to_unsigned( 176, 8)),
10 => std_logic_vector(to_unsigned( 75, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 255, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 52, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 85 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 116, 8)),
2 => std_logic_vector(to_unsigned( 216, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 74, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 241, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 163, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 169, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 86 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 14, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 66, 8)),
5 => std_logic_vector(to_unsigned( 88, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 150, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 87 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 76, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 31, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 21, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 25, 8)),
10 => std_logic_vector(to_unsigned( 100, 8)),
11 => std_logic_vector(to_unsigned( 40, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 16, 8)),
16 => std_logic_vector(to_unsigned( 214, 8)),
17 => std_logic_vector(to_unsigned( 52, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 88 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 0, 8)),
4 => std_logic_vector(to_unsigned( 77, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 198, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 188, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 155, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 188, 8)),
18 => std_logic_vector(to_unsigned( 106, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 89 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 64, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 239, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 208, 8)),
10 => std_logic_vector(to_unsigned( 244, 8)),
11 => std_logic_vector(to_unsigned( 247, 8)),
12 => std_logic_vector(to_unsigned( 66, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 163, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 90 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 157, 8)),
3 => std_logic_vector(to_unsigned( 131, 8)),
4 => std_logic_vector(to_unsigned( 187, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 165, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 59, 8)),
15 => std_logic_vector(to_unsigned( 212, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 91 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 227, 8)),
3 => std_logic_vector(to_unsigned( 186, 8)),
4 => std_logic_vector(to_unsigned( 223, 8)),
5 => std_logic_vector(to_unsigned( 235, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 103, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 72, 8)),
10 => std_logic_vector(to_unsigned( 52, 8)),
11 => std_logic_vector(to_unsigned( 199, 8)),
12 => std_logic_vector(to_unsigned( 210, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 92 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 108, 8)),
5 => std_logic_vector(to_unsigned( 43, 8)),
6 => std_logic_vector(to_unsigned( 232, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 216, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 1, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 74, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 33, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 93 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 23, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 189, 8)),
6 => std_logic_vector(to_unsigned( 172, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 137, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 145, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 48, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 94 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 229, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 29, 8)),
5 => std_logic_vector(to_unsigned( 42, 8)),
6 => std_logic_vector(to_unsigned( 45, 8)),
7 => std_logic_vector(to_unsigned( 78, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 1, 8)),
11 => std_logic_vector(to_unsigned( 92, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 95 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 211, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 244, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 212, 8)),
8 => std_logic_vector(to_unsigned( 54, 8)),
9 => std_logic_vector(to_unsigned( 118, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 198, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 191, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 96 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 83, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 113, 8)),
4 => std_logic_vector(to_unsigned( 12, 8)),
5 => std_logic_vector(to_unsigned( 142, 8)),
6 => std_logic_vector(to_unsigned( 142, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 172, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 209, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 97 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 27, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 34, 8)),
4 => std_logic_vector(to_unsigned( 241, 8)),
5 => std_logic_vector(to_unsigned( 72, 8)),
6 => std_logic_vector(to_unsigned( 33, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 38, 8)),
12 => std_logic_vector(to_unsigned( 225, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 230, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 233, 8)),
17 => std_logic_vector(to_unsigned( 55, 8)),
18 => std_logic_vector(to_unsigned( 212, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 98 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 136, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 170, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 229, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 118, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 99 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 215, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 215, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 115, 8)),
7 => std_logic_vector(to_unsigned( 148, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 138, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 192, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 58, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 100 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 9, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 88, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 172, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 39, 8)),
10 => std_logic_vector(to_unsigned( 16, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100110
elsif count = 101 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 199, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 207, 8)),
6 => std_logic_vector(to_unsigned( 204, 8)),
7 => std_logic_vector(to_unsigned( 207, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 3, 8)),
11 => std_logic_vector(to_unsigned( 76, 8)),
12 => std_logic_vector(to_unsigned( 90, 8)),
13 => std_logic_vector(to_unsigned( 14, 8)),
14 => std_logic_vector(to_unsigned( 239, 8)),
15 => std_logic_vector(to_unsigned( 152, 8)),
16 => std_logic_vector(to_unsigned( 11, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 56, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001011
elsif count = 102 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 166, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 89, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 203, 8)),
13 => std_logic_vector(to_unsigned( 60, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 103 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 61, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 157, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 238, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 226, 8)),
14 => std_logic_vector(to_unsigned( 85, 8)),
15 => std_logic_vector(to_unsigned( 16, 8)),
16 => std_logic_vector(to_unsigned( 185, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 104 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 214, 8)),
10 => std_logic_vector(to_unsigned( 87, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 248, 8)),
14 => std_logic_vector(to_unsigned( 163, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 81, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 105 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 4, 8)),
3 => std_logic_vector(to_unsigned( 209, 8)),
4 => std_logic_vector(to_unsigned( 26, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 168, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 165, 8)),
11 => std_logic_vector(to_unsigned( 11, 8)),
12 => std_logic_vector(to_unsigned( 85, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 106 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 239, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 27, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 205, 8)),
12 => std_logic_vector(to_unsigned( 48, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 46, 8)),
16 => std_logic_vector(to_unsigned( 238, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111100
elsif count = 107 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 35, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 155, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 173, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 230, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 27, 8)),
17 => std_logic_vector(to_unsigned( 75, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 108 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 28, 8)),
4 => std_logic_vector(to_unsigned( 178, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 38, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 131, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 108, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 109 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 79, 8)),
2 => std_logic_vector(to_unsigned( 191, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 254, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 235, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 101, 8)),
12 => std_logic_vector(to_unsigned( 223, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 241, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 110 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 197, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 177, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 203, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 50, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 111 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 78, 8)),
2 => std_logic_vector(to_unsigned( 192, 8)),
3 => std_logic_vector(to_unsigned( 27, 8)),
4 => std_logic_vector(to_unsigned( 47, 8)),
5 => std_logic_vector(to_unsigned( 13, 8)),
6 => std_logic_vector(to_unsigned( 87, 8)),
7 => std_logic_vector(to_unsigned( 64, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 231, 8)),
10 => std_logic_vector(to_unsigned( 6, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 69, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 56, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 112 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 203, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 63, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 216, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 42, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 60, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 8, 8)),
14 => std_logic_vector(to_unsigned( 75, 8)),
15 => std_logic_vector(to_unsigned( 204, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 113 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 144, 8)),
3 => std_logic_vector(to_unsigned( 254, 8)),
4 => std_logic_vector(to_unsigned( 193, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 180, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 2, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 239, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 114 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 89, 8)),
4 => std_logic_vector(to_unsigned( 117, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 94, 8)),
11 => std_logic_vector(to_unsigned( 78, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 220, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 11, 8)),
16 => std_logic_vector(to_unsigned( 213, 8)),
17 => std_logic_vector(to_unsigned( 81, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 115 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 87, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 4, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 15, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 187, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 29, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 116 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 75, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 240, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 83, 8)),
7 => std_logic_vector(to_unsigned( 237, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 115, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 102, 8)),
17 => std_logic_vector(to_unsigned( 206, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 117 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 197, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 184, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 139, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 63, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 105, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 118 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 19, 8)),
4 => std_logic_vector(to_unsigned( 64, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 63, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 141, 8)),
14 => std_logic_vector(to_unsigned( 145, 8)),
15 => std_logic_vector(to_unsigned( 193, 8)),
16 => std_logic_vector(to_unsigned( 79, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111100
elsif count = 119 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 75, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 226, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 193, 8)),
9 => std_logic_vector(to_unsigned( 114, 8)),
10 => std_logic_vector(to_unsigned( 107, 8)),
11 => std_logic_vector(to_unsigned( 150, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 26, 8)),
14 => std_logic_vector(to_unsigned( 85, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 81, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 120 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 23, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 197, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 184, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 252, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 177, 8)),
15 => std_logic_vector(to_unsigned( 200, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 181, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 121 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 47, 8)),
4 => std_logic_vector(to_unsigned( 218, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 170, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 173, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 71, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 214, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 122 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 205, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 200, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 117, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 197, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 207, 8)),
11 => std_logic_vector(to_unsigned( 240, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 239, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 185, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 123 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 35, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 41, 8)),
8 => std_logic_vector(to_unsigned( 82, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 41, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 197, 8)),
14 => std_logic_vector(to_unsigned( 140, 8)),
15 => std_logic_vector(to_unsigned( 235, 8)),
16 => std_logic_vector(to_unsigned( 195, 8)),
17 => std_logic_vector(to_unsigned( 41, 8)),
18 => std_logic_vector(to_unsigned( 41, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 124 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 196, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 173, 8)),
7 => std_logic_vector(to_unsigned( 87, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 146, 8)),
10 => std_logic_vector(to_unsigned( 244, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 125 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 129, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 243, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 116, 8)),
13 => std_logic_vector(to_unsigned( 66, 8)),
14 => std_logic_vector(to_unsigned( 80, 8)),
15 => std_logic_vector(to_unsigned( 98, 8)),
16 => std_logic_vector(to_unsigned( 162, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 126 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 131, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 183, 8)),
6 => std_logic_vector(to_unsigned( 2, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 63, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 40, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 127 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 205, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 176, 8)),
8 => std_logic_vector(to_unsigned( 92, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 77, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 36, 8)),
13 => std_logic_vector(to_unsigned( 242, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 27, 8)),
17 => std_logic_vector(to_unsigned( 189, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 128 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 43, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 49, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 162, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 13, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 129 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 30, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 211, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 53, 8)),
7 => std_logic_vector(to_unsigned( 39, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 249, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 57, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 36, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 130 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 70, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 201, 8)),
4 => std_logic_vector(to_unsigned( 219, 8)),
5 => std_logic_vector(to_unsigned( 227, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 85, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 107, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 84, 8)),
13 => std_logic_vector(to_unsigned( 186, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 182, 8)),
16 => std_logic_vector(to_unsigned( 59, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 131 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 20, 8)),
2 => std_logic_vector(to_unsigned( 240, 8)),
3 => std_logic_vector(to_unsigned( 36, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 184, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 230, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 245, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 119, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 132 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 33, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 111, 8)),
10 => std_logic_vector(to_unsigned( 122, 8)),
11 => std_logic_vector(to_unsigned( 147, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 15, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 133 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 91, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 150, 8)),
8 => std_logic_vector(to_unsigned( 89, 8)),
9 => std_logic_vector(to_unsigned( 56, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 230, 8)),
14 => std_logic_vector(to_unsigned( 12, 8)),
15 => std_logic_vector(to_unsigned( 191, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 134 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 27, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 221, 8)),
4 => std_logic_vector(to_unsigned( 203, 8)),
5 => std_logic_vector(to_unsigned( 170, 8)),
6 => std_logic_vector(to_unsigned( 240, 8)),
7 => std_logic_vector(to_unsigned( 78, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 255, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 219, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 173, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 211, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 135 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 210, 8)),
10 => std_logic_vector(to_unsigned( 234, 8)),
11 => std_logic_vector(to_unsigned( 70, 8)),
12 => std_logic_vector(to_unsigned( 95, 8)),
13 => std_logic_vector(to_unsigned( 226, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 216, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001100
elsif count = 136 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 45, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 203, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 229, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 5, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 175, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 182, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 137 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 88, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 246, 8)),
10 => std_logic_vector(to_unsigned( 159, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 80, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 10, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00100111
elsif count = 138 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 226, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 3, 8)),
13 => std_logic_vector(to_unsigned( 138, 8)),
14 => std_logic_vector(to_unsigned( 248, 8)),
15 => std_logic_vector(to_unsigned( 211, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 182, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 139 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 22, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 12, 8)),
5 => std_logic_vector(to_unsigned( 82, 8)),
6 => std_logic_vector(to_unsigned( 112, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 138, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 140 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 144, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 105, 8)),
5 => std_logic_vector(to_unsigned( 20, 8)),
6 => std_logic_vector(to_unsigned( 11, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 178, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 141 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 17, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 18, 8)),
9 => std_logic_vector(to_unsigned( 186, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 142 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 214, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 16, 8)),
4 => std_logic_vector(to_unsigned( 73, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 190, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 209, 8)),
15 => std_logic_vector(to_unsigned( 27, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 143 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 163, 8)),
2 => std_logic_vector(to_unsigned( 38, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 170, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 87, 8)),
11 => std_logic_vector(to_unsigned( 199, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 144 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 185, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 182, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 54, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 79, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 145 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 241, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 16, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 119, 8)),
11 => std_logic_vector(to_unsigned( 7, 8)),
12 => std_logic_vector(to_unsigned( 233, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 190, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011010
elsif count = 146 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 230, 8)),
2 => std_logic_vector(to_unsigned( 249, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 92, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 43, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 243, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 34, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 68, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 61, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 147 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 184, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 13, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 211, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 91, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 148 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 195, 8)),
2 => std_logic_vector(to_unsigned( 61, 8)),
3 => std_logic_vector(to_unsigned( 204, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 215, 8)),
6 => std_logic_vector(to_unsigned( 14, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 234, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 111, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 232, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 149 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 158, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 195, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 31, 8)),
11 => std_logic_vector(to_unsigned( 41, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 59, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 150 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 54, 8)),
2 => std_logic_vector(to_unsigned( 178, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 233, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 87, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 74, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010110
elsif count = 151 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 99, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 179, 8)),
6 => std_logic_vector(to_unsigned( 87, 8)),
7 => std_logic_vector(to_unsigned( 27, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 152 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 19, 8)),
3 => std_logic_vector(to_unsigned( 129, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 227, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 77, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 37, 8)),
15 => std_logic_vector(to_unsigned( 55, 8)),
16 => std_logic_vector(to_unsigned( 119, 8)),
17 => std_logic_vector(to_unsigned( 75, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100010
elsif count = 153 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 66, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 73, 8)),
4 => std_logic_vector(to_unsigned( 242, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 53, 8)),
8 => std_logic_vector(to_unsigned( 189, 8)),
9 => std_logic_vector(to_unsigned( 96, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 154 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 42, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 100, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 101, 8)),
6 => std_logic_vector(to_unsigned( 208, 8)),
7 => std_logic_vector(to_unsigned( 71, 8)),
8 => std_logic_vector(to_unsigned( 178, 8)),
9 => std_logic_vector(to_unsigned( 132, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 74, 8)),
14 => std_logic_vector(to_unsigned( 151, 8)),
15 => std_logic_vector(to_unsigned( 10, 8)),
16 => std_logic_vector(to_unsigned( 102, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 155 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 45, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 40, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 160, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 245, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 75, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 156 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 48, 8)),
6 => std_logic_vector(to_unsigned( 225, 8)),
7 => std_logic_vector(to_unsigned( 77, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 39, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 12, 8)),
12 => std_logic_vector(to_unsigned( 193, 8)),
13 => std_logic_vector(to_unsigned( 10, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 185, 8)),
16 => std_logic_vector(to_unsigned( 35, 8)),
17 => std_logic_vector(to_unsigned( 46, 8)),
18 => std_logic_vector(to_unsigned( 190, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 157 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 3, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 28, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 12, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 28, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 48, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 40, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 158 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 58, 8)),
7 => std_logic_vector(to_unsigned( 85, 8)),
8 => std_logic_vector(to_unsigned( 75, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 79, 8)),
14 => std_logic_vector(to_unsigned( 69, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 11, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 159 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 228, 8)),
2 => std_logic_vector(to_unsigned( 160, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 2, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 54, 8)),
12 => std_logic_vector(to_unsigned( 78, 8)),
13 => std_logic_vector(to_unsigned( 141, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 160 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 88, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 210, 8)),
8 => std_logic_vector(to_unsigned( 22, 8)),
9 => std_logic_vector(to_unsigned( 82, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 48, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 161 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 219, 8)),
4 => std_logic_vector(to_unsigned( 184, 8)),
5 => std_logic_vector(to_unsigned( 211, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 203, 8)),
8 => std_logic_vector(to_unsigned( 230, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 227, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 179, 8)),
14 => std_logic_vector(to_unsigned( 21, 8)),
15 => std_logic_vector(to_unsigned( 229, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 200, 8)),
18 => std_logic_vector(to_unsigned( 199, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 162 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 14, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 162, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 239, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101100
elsif count = 163 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 136, 8)),
2 => std_logic_vector(to_unsigned( 171, 8)),
3 => std_logic_vector(to_unsigned( 76, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 119, 8)),
11 => std_logic_vector(to_unsigned( 38, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 220, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 164 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 36, 8)),
5 => std_logic_vector(to_unsigned( 119, 8)),
6 => std_logic_vector(to_unsigned( 20, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 30, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 77, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 41, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 165 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 238, 8)),
2 => std_logic_vector(to_unsigned( 23, 8)),
3 => std_logic_vector(to_unsigned( 15, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 194, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 112, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 166 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 82, 8)),
3 => std_logic_vector(to_unsigned( 109, 8)),
4 => std_logic_vector(to_unsigned( 6, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 87, 8)),
12 => std_logic_vector(to_unsigned( 68, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 20, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 5, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 47, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 167 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 171, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 106, 8)),
5 => std_logic_vector(to_unsigned( 47, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 3, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 217, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 140, 8)),
13 => std_logic_vector(to_unsigned( 73, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 168 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 236, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 20, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 222, 8)),
7 => std_logic_vector(to_unsigned( 244, 8)),
8 => std_logic_vector(to_unsigned( 77, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 141, 8)),
14 => std_logic_vector(to_unsigned( 226, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 123, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 169 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 229, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 182, 8)),
7 => std_logic_vector(to_unsigned( 244, 8)),
8 => std_logic_vector(to_unsigned( 24, 8)),
9 => std_logic_vector(to_unsigned( 134, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 217, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 131, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 170 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 26, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 227, 8)),
8 => std_logic_vector(to_unsigned( 193, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 12, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 171 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 13, 8)),
5 => std_logic_vector(to_unsigned( 181, 8)),
6 => std_logic_vector(to_unsigned( 25, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 109, 8)),
9 => std_logic_vector(to_unsigned( 217, 8)),
10 => std_logic_vector(to_unsigned( 211, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 23, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 172 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 31, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 31, 8)),
4 => std_logic_vector(to_unsigned( 74, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 89, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 42, 8)),
14 => std_logic_vector(to_unsigned( 218, 8)),
15 => std_logic_vector(to_unsigned( 58, 8)),
16 => std_logic_vector(to_unsigned( 174, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 173 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 197, 8)),
2 => std_logic_vector(to_unsigned( 182, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 62, 8)),
5 => std_logic_vector(to_unsigned( 248, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 202, 8)),
8 => std_logic_vector(to_unsigned( 140, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 221, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 151, 8)),
13 => std_logic_vector(to_unsigned( 135, 8)),
14 => std_logic_vector(to_unsigned( 216, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 174 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 63, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 242, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 250, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 39, 8)),
16 => std_logic_vector(to_unsigned( 235, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00010111
elsif count = 175 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 145, 8)),
3 => std_logic_vector(to_unsigned( 8, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 251, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 23, 8)),
11 => std_logic_vector(to_unsigned( 150, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 54, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 176 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 239, 8)),
2 => std_logic_vector(to_unsigned( 155, 8)),
3 => std_logic_vector(to_unsigned( 210, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 209, 8)),
7 => std_logic_vector(to_unsigned( 147, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 246, 8)),
10 => std_logic_vector(to_unsigned( 239, 8)),
11 => std_logic_vector(to_unsigned( 183, 8)),
12 => std_logic_vector(to_unsigned( 249, 8)),
13 => std_logic_vector(to_unsigned( 157, 8)),
14 => std_logic_vector(to_unsigned( 179, 8)),
15 => std_logic_vector(to_unsigned( 143, 8)),
16 => std_logic_vector(to_unsigned( 178, 8)),
17 => std_logic_vector(to_unsigned( 188, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 177 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 26, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 89, 8)),
8 => std_logic_vector(to_unsigned( 220, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 178 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 69, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 38, 8)),
5 => std_logic_vector(to_unsigned( 190, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 225, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 68, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 216, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 184, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 179 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 209, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 254, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 53, 8)),
13 => std_logic_vector(to_unsigned( 152, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 231, 8)),
16 => std_logic_vector(to_unsigned( 161, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00010111
elsif count = 180 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 71, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 209, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 15, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 245, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 90, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 128, 8)),
15 => std_logic_vector(to_unsigned( 72, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 181 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 241, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 83, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 51, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 226, 8)),
12 => std_logic_vector(to_unsigned( 208, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 81, 8)),
16 => std_logic_vector(to_unsigned( 202, 8)),
17 => std_logic_vector(to_unsigned( 73, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 182 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 207, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 162, 8)),
4 => std_logic_vector(to_unsigned( 224, 8)),
5 => std_logic_vector(to_unsigned( 235, 8)),
6 => std_logic_vector(to_unsigned( 44, 8)),
7 => std_logic_vector(to_unsigned( 177, 8)),
8 => std_logic_vector(to_unsigned( 253, 8)),
9 => std_logic_vector(to_unsigned( 216, 8)),
10 => std_logic_vector(to_unsigned( 124, 8)),
11 => std_logic_vector(to_unsigned( 161, 8)),
12 => std_logic_vector(to_unsigned( 151, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 131, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 183 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 197, 8)),
2 => std_logic_vector(to_unsigned( 250, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 32, 8)),
7 => std_logic_vector(to_unsigned( 108, 8)),
8 => std_logic_vector(to_unsigned( 45, 8)),
9 => std_logic_vector(to_unsigned( 63, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 18, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 52, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 48, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 61, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 184 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 13, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 112, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 123, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 32, 8)),
9 => std_logic_vector(to_unsigned( 45, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 13, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 240, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 185 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 216, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 254, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 13, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 33, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 46, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 186 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 82, 8)),
9 => std_logic_vector(to_unsigned( 138, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 45, 8)),
12 => std_logic_vector(to_unsigned( 249, 8)),
13 => std_logic_vector(to_unsigned( 211, 8)),
14 => std_logic_vector(to_unsigned( 198, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 187 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 243, 8)),
2 => std_logic_vector(to_unsigned( 234, 8)),
3 => std_logic_vector(to_unsigned( 38, 8)),
4 => std_logic_vector(to_unsigned( 238, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 202, 8)),
8 => std_logic_vector(to_unsigned( 56, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 101, 8)),
12 => std_logic_vector(to_unsigned( 75, 8)),
13 => std_logic_vector(to_unsigned( 152, 8)),
14 => std_logic_vector(to_unsigned( 126, 8)),
15 => std_logic_vector(to_unsigned( 218, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 188 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 147, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 43, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 58, 8)),
9 => std_logic_vector(to_unsigned( 214, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 63, 8)),
12 => std_logic_vector(to_unsigned( 98, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 13, 8)),
16 => std_logic_vector(to_unsigned( 251, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 189 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 204, 8)),
2 => std_logic_vector(to_unsigned( 156, 8)),
3 => std_logic_vector(to_unsigned( 193, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 132, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 210, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 190 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 36, 8)),
3 => std_logic_vector(to_unsigned( 75, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 71, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 5, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 167, 8)),
12 => std_logic_vector(to_unsigned( 58, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 227, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 37, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 191 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 94, 8)),
3 => std_logic_vector(to_unsigned( 150, 8)),
4 => std_logic_vector(to_unsigned( 90, 8)),
5 => std_logic_vector(to_unsigned( 26, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 243, 8)),
8 => std_logic_vector(to_unsigned( 81, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 169, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 131, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 192 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 14, 8)),
6 => std_logic_vector(to_unsigned( 206, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 198, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 225, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 245, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 193 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 199, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 7, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 253, 8)),
9 => std_logic_vector(to_unsigned( 215, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 203, 8)),
12 => std_logic_vector(to_unsigned( 62, 8)),
13 => std_logic_vector(to_unsigned( 98, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 197, 8)),
16 => std_logic_vector(to_unsigned( 58, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 194 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 26, 8)),
4 => std_logic_vector(to_unsigned( 20, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 232, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 249, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100100
elsif count = 195 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 77, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 18, 8)),
10 => std_logic_vector(to_unsigned( 254, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 41, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 100, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 196 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 195, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 1, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 219, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 136, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 152, 8)),
15 => std_logic_vector(to_unsigned( 213, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 197 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 11, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 209, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 214, 8)),
9 => std_logic_vector(to_unsigned( 136, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 165, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 183, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 198 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 249, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 195, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 228, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 181, 8)),
12 => std_logic_vector(to_unsigned( 221, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 58, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 199 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 190, 8)),
2 => std_logic_vector(to_unsigned( 34, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 50, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 76, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 12, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 59, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 200 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 56, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 112, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 41, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 37, 8)),
15 => std_logic_vector(to_unsigned( 18, 8)),
16 => std_logic_vector(to_unsigned( 252, 8)),
17 => std_logic_vector(to_unsigned( 75, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110110
elsif count = 201 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 28, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 66, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 239, 8)),
12 => std_logic_vector(to_unsigned( 245, 8)),
13 => std_logic_vector(to_unsigned( 190, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 202 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 30, 8)),
3 => std_logic_vector(to_unsigned( 30, 8)),
4 => std_logic_vector(to_unsigned( 29, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 245, 8)),
8 => std_logic_vector(to_unsigned( 243, 8)),
9 => std_logic_vector(to_unsigned( 4, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 215, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 225, 8)),
17 => std_logic_vector(to_unsigned( 41, 8)),
18 => std_logic_vector(to_unsigned( 58, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00010111
elsif count = 203 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 98, 8)),
4 => std_logic_vector(to_unsigned( 90, 8)),
5 => std_logic_vector(to_unsigned( 77, 8)),
6 => std_logic_vector(to_unsigned( 224, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 127, 8)),
9 => std_logic_vector(to_unsigned( 34, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 160, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 173, 8)),
16 => std_logic_vector(to_unsigned( 145, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 204 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 157, 8)),
4 => std_logic_vector(to_unsigned( 26, 8)),
5 => std_logic_vector(to_unsigned( 173, 8)),
6 => std_logic_vector(to_unsigned( 10, 8)),
7 => std_logic_vector(to_unsigned( 213, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 42, 8)),
10 => std_logic_vector(to_unsigned( 23, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 13, 8)),
13 => std_logic_vector(to_unsigned( 228, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 234, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 205 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 238, 8)),
3 => std_logic_vector(to_unsigned( 80, 8)),
4 => std_logic_vector(to_unsigned( 247, 8)),
5 => std_logic_vector(to_unsigned( 14, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 228, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 180, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 254, 8)),
15 => std_logic_vector(to_unsigned( 247, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 190, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 206 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 181, 8)),
8 => std_logic_vector(to_unsigned( 182, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 95, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 207 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 211, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 0, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 7, 8)),
8 => std_logic_vector(to_unsigned( 182, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 78, 8)),
18 => std_logic_vector(to_unsigned( 183, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 208 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 186, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 159, 8)),
4 => std_logic_vector(to_unsigned( 223, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 245, 8)),
8 => std_logic_vector(to_unsigned( 89, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 235, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 213, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 205, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 209 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 141, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 244, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 245, 8)),
8 => std_logic_vector(to_unsigned( 18, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 118, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 210 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 169, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 82, 8)),
9 => std_logic_vector(to_unsigned( 218, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 211 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 95, 8)),
2 => std_logic_vector(to_unsigned( 224, 8)),
3 => std_logic_vector(to_unsigned( 178, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 141, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 110, 8)),
10 => std_logic_vector(to_unsigned( 239, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 40, 8)),
13 => std_logic_vector(to_unsigned( 73, 8)),
14 => std_logic_vector(to_unsigned( 202, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010111
elsif count = 212 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 71, 8)),
2 => std_logic_vector(to_unsigned( 254, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 20, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 184, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 68, 8)),
13 => std_logic_vector(to_unsigned( 69, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 213 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 31, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 36, 8)),
6 => std_logic_vector(to_unsigned( 152, 8)),
7 => std_logic_vector(to_unsigned( 53, 8)),
8 => std_logic_vector(to_unsigned( 197, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 183, 8)),
11 => std_logic_vector(to_unsigned( 38, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 10, 8)),
14 => std_logic_vector(to_unsigned( 186, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 75, 8)),
17 => std_logic_vector(to_unsigned( 37, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 214 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 2, 8)),
2 => std_logic_vector(to_unsigned( 6, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 134, 8)),
7 => std_logic_vector(to_unsigned( 14, 8)),
8 => std_logic_vector(to_unsigned( 106, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 156, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 40, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 215 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 242, 8)),
4 => std_logic_vector(to_unsigned( 183, 8)),
5 => std_logic_vector(to_unsigned( 100, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 234, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 66, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 87, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 156, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 79, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 216 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 187, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 5, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 212, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 3, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 210, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 184, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 217 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 215, 8)),
3 => std_logic_vector(to_unsigned( 213, 8)),
4 => std_logic_vector(to_unsigned( 244, 8)),
5 => std_logic_vector(to_unsigned( 7, 8)),
6 => std_logic_vector(to_unsigned( 255, 8)),
7 => std_logic_vector(to_unsigned( 216, 8)),
8 => std_logic_vector(to_unsigned( 253, 8)),
9 => std_logic_vector(to_unsigned( 84, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 218 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 162, 8)),
2 => std_logic_vector(to_unsigned( 144, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 41, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 215, 8)),
8 => std_logic_vector(to_unsigned( 48, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 35, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 79, 8)),
13 => std_logic_vector(to_unsigned( 222, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 53, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 219 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 34, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 158, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 238, 8)),
8 => std_logic_vector(to_unsigned( 226, 8)),
9 => std_logic_vector(to_unsigned( 30, 8)),
10 => std_logic_vector(to_unsigned( 74, 8)),
11 => std_logic_vector(to_unsigned( 57, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 1, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 58, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010110
elsif count = 220 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 254, 8)),
5 => std_logic_vector(to_unsigned( 216, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 163, 8)),
14 => std_logic_vector(to_unsigned( 214, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 191, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 221 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 202, 8)),
5 => std_logic_vector(to_unsigned( 109, 8)),
6 => std_logic_vector(to_unsigned( 189, 8)),
7 => std_logic_vector(to_unsigned( 214, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 180, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 126, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 207, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 222 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 230, 8)),
3 => std_logic_vector(to_unsigned( 25, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 75, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 107, 8)),
11 => std_logic_vector(to_unsigned( 132, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 144, 8)),
15 => std_logic_vector(to_unsigned( 54, 8)),
16 => std_logic_vector(to_unsigned( 190, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 223 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 177, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 247, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 107, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 204, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 178, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 224 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 72, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 224, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 3, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 234, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001011
elsif count = 225 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 20, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 32, 8)),
4 => std_logic_vector(to_unsigned( 250, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 23, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 77, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 48, 8)),
13 => std_logic_vector(to_unsigned( 34, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 56, 8)),
16 => std_logic_vector(to_unsigned( 132, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 226 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 205, 8)),
3 => std_logic_vector(to_unsigned( 75, 8)),
4 => std_logic_vector(to_unsigned( 209, 8)),
5 => std_logic_vector(to_unsigned( 103, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 184, 8)),
8 => std_logic_vector(to_unsigned( 211, 8)),
9 => std_logic_vector(to_unsigned( 202, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 210, 8)),
12 => std_logic_vector(to_unsigned( 191, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 168, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 227 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 36, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 103, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 28, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 204, 8)),
13 => std_logic_vector(to_unsigned( 71, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 228, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 228 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 47, 8)),
2 => std_logic_vector(to_unsigned( 197, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 16, 8)),
5 => std_logic_vector(to_unsigned( 116, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 22, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 232, 8)),
10 => std_logic_vector(to_unsigned( 23, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 39, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 51, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 229 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 251, 8)),
3 => std_logic_vector(to_unsigned( 213, 8)),
4 => std_logic_vector(to_unsigned( 28, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 127, 8)),
16 => std_logic_vector(to_unsigned( 215, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 230 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 210, 8)),
3 => std_logic_vector(to_unsigned( 169, 8)),
4 => std_logic_vector(to_unsigned( 193, 8)),
5 => std_logic_vector(to_unsigned( 82, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 20, 8)),
8 => std_logic_vector(to_unsigned( 206, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 170, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 231 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 81, 8)),
4 => std_logic_vector(to_unsigned( 234, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 131, 8)),
12 => std_logic_vector(to_unsigned( 204, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 252, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011101
elsif count = 232 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 46, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 197, 8)),
6 => std_logic_vector(to_unsigned( 231, 8)),
7 => std_logic_vector(to_unsigned( 161, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 109, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 45, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 74, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110000
elsif count = 233 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 182, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 192, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 189, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 182, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 234 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 225, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 48, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 77, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 34, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 55, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 50, 8)),
16 => std_logic_vector(to_unsigned( 235, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101110
elsif count = 235 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 129, 8)),
2 => std_logic_vector(to_unsigned( 238, 8)),
3 => std_logic_vector(to_unsigned( 49, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 189, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 45, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 59, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001100
elsif count = 236 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 246, 8)),
2 => std_logic_vector(to_unsigned( 34, 8)),
3 => std_logic_vector(to_unsigned( 70, 8)),
4 => std_logic_vector(to_unsigned( 245, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 34, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 35, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 27, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 81, 8)),
13 => std_logic_vector(to_unsigned( 18, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 252, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111100
elsif count = 237 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 32, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 28, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 11, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 196, 8)),
11 => std_logic_vector(to_unsigned( 24, 8)),
12 => std_logic_vector(to_unsigned( 180, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 58, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 238 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 64, 8)),
3 => std_logic_vector(to_unsigned( 140, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 135, 8)),
8 => std_logic_vector(to_unsigned( 49, 8)),
9 => std_logic_vector(to_unsigned( 39, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 129, 8)),
12 => std_logic_vector(to_unsigned( 179, 8)),
13 => std_logic_vector(to_unsigned( 100, 8)),
14 => std_logic_vector(to_unsigned( 73, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 239 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 212, 8)),
3 => std_logic_vector(to_unsigned( 240, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 40, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 67, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 247, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 26, 8)),
16 => std_logic_vector(to_unsigned( 13, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 240 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 220, 8)),
3 => std_logic_vector(to_unsigned( 99, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 243, 8)),
6 => std_logic_vector(to_unsigned( 212, 8)),
7 => std_logic_vector(to_unsigned( 89, 8)),
8 => std_logic_vector(to_unsigned( 106, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 24, 8)),
11 => std_logic_vector(to_unsigned( 63, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 136, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 241 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 13, 8)),
3 => std_logic_vector(to_unsigned( 84, 8)),
4 => std_logic_vector(to_unsigned( 177, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 30, 8)),
7 => std_logic_vector(to_unsigned( 223, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 172, 8)),
12 => std_logic_vector(to_unsigned( 225, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 172, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 231, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110010
elsif count = 242 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 217, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 90, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 218, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 202, 8)),
8 => std_logic_vector(to_unsigned( 253, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 215, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 39, 8)),
16 => std_logic_vector(to_unsigned( 202, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 243 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 233, 8)),
2 => std_logic_vector(to_unsigned( 220, 8)),
3 => std_logic_vector(to_unsigned( 27, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 11, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 206, 8)),
10 => std_logic_vector(to_unsigned( 178, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 244 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 55, 8)),
3 => std_logic_vector(to_unsigned( 201, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 46, 8)),
6 => std_logic_vector(to_unsigned( 23, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 69, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 255, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 61, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 245 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 221, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 81, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 246 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 38, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 89, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 70, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 16, 8)),
15 => std_logic_vector(to_unsigned( 8, 8)),
16 => std_logic_vector(to_unsigned( 217, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 247 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 251, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 237, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 224, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 73, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 248 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 6, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 44, 8)),
11 => std_logic_vector(to_unsigned( 83, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 79, 8)),
14 => std_logic_vector(to_unsigned( 119, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 249 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 71, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 219, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 214, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 216, 8)),
16 => std_logic_vector(to_unsigned( 192, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 201, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 250 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 220, 8)),
2 => std_logic_vector(to_unsigned( 246, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 34, 8)),
5 => std_logic_vector(to_unsigned( 93, 8)),
6 => std_logic_vector(to_unsigned( 117, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 173, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 45, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 34, 8)),
15 => std_logic_vector(to_unsigned( 5, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 251 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 83, 8)),
4 => std_logic_vector(to_unsigned( 192, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 28, 8)),
7 => std_logic_vector(to_unsigned( 116, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 7, 8)),
10 => std_logic_vector(to_unsigned( 89, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 96, 8)),
13 => std_logic_vector(to_unsigned( 222, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 131, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 252 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 36, 8)),
4 => std_logic_vector(to_unsigned( 177, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 37, 8)),
13 => std_logic_vector(to_unsigned( 95, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 193, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 253 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 185, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 222, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 86, 8)),
10 => std_logic_vector(to_unsigned( 248, 8)),
11 => std_logic_vector(to_unsigned( 228, 8)),
12 => std_logic_vector(to_unsigned( 140, 8)),
13 => std_logic_vector(to_unsigned( 157, 8)),
14 => std_logic_vector(to_unsigned( 215, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 254 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 170, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 32, 8)),
4 => std_logic_vector(to_unsigned( 241, 8)),
5 => std_logic_vector(to_unsigned( 77, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 132, 8)),
8 => std_logic_vector(to_unsigned( 30, 8)),
9 => std_logic_vector(to_unsigned( 77, 8)),
10 => std_logic_vector(to_unsigned( 245, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 63, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 255 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 214, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 156, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 1, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 256 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 250, 8)),
2 => std_logic_vector(to_unsigned( 51, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 64, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 252, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 224, 8)),
12 => std_logic_vector(to_unsigned( 37, 8)),
13 => std_logic_vector(to_unsigned( 217, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 257 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 220, 8)),
3 => std_logic_vector(to_unsigned( 80, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 53, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 155, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 130, 8)),
15 => std_logic_vector(to_unsigned( 185, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101110
elsif count = 258 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 29, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 140, 8)),
4 => std_logic_vector(to_unsigned( 72, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 226, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 190, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 163, 8)),
14 => std_logic_vector(to_unsigned( 45, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 51, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 259 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 230, 8)),
8 => std_logic_vector(to_unsigned( 61, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 76, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 179, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011001
elsif count = 260 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 14, 8)),
2 => std_logic_vector(to_unsigned( 42, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 25, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 167, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 52, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100010
elsif count = 261 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 36, 8)),
3 => std_logic_vector(to_unsigned( 224, 8)),
4 => std_logic_vector(to_unsigned( 59, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 50, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 86, 8)),
9 => std_logic_vector(to_unsigned( 215, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 200, 8)),
12 => std_logic_vector(to_unsigned( 35, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 50, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 262 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 29, 8)),
5 => std_logic_vector(to_unsigned( 219, 8)),
6 => std_logic_vector(to_unsigned( 224, 8)),
7 => std_logic_vector(to_unsigned( 211, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 223, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 152, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 164, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 118, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 263 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 194, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 28, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 216, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 264 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 180, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 242, 8)),
8 => std_logic_vector(to_unsigned( 112, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 6, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 136, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 185, 8)),
16 => std_logic_vector(to_unsigned( 173, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 265 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 45, 8)),
3 => std_logic_vector(to_unsigned( 227, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 247, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 237, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 220, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 24, 8)),
16 => std_logic_vector(to_unsigned( 19, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 266 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 12, 8)),
2 => std_logic_vector(to_unsigned( 52, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 208, 8)),
5 => std_logic_vector(to_unsigned( 148, 8)),
6 => std_logic_vector(to_unsigned( 24, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 179, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 147, 8)),
12 => std_logic_vector(to_unsigned( 27, 8)),
13 => std_logic_vector(to_unsigned( 197, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 133, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 267 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 207, 8)),
5 => std_logic_vector(to_unsigned( 100, 8)),
6 => std_logic_vector(to_unsigned( 227, 8)),
7 => std_logic_vector(to_unsigned( 24, 8)),
8 => std_logic_vector(to_unsigned( 220, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 224, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 205, 8)),
15 => std_logic_vector(to_unsigned( 245, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 268 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 242, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 162, 8)),
4 => std_logic_vector(to_unsigned( 41, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 21, 8)),
8 => std_logic_vector(to_unsigned( 155, 8)),
9 => std_logic_vector(to_unsigned( 85, 8)),
10 => std_logic_vector(to_unsigned( 116, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 41, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 269 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 61, 8)),
3 => std_logic_vector(to_unsigned( 200, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 244, 8)),
10 => std_logic_vector(to_unsigned( 251, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 270 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 2, 8)),
2 => std_logic_vector(to_unsigned( 207, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 197, 8)),
6 => std_logic_vector(to_unsigned( 114, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 89, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 30, 8)),
13 => std_logic_vector(to_unsigned( 150, 8)),
14 => std_logic_vector(to_unsigned( 4, 8)),
15 => std_logic_vector(to_unsigned( 99, 8)),
16 => std_logic_vector(to_unsigned( 12, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 271 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 143, 8)),
3 => std_logic_vector(to_unsigned( 10, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 1, 8)),
6 => std_logic_vector(to_unsigned( 28, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 90, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 74, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 77, 8)),
15 => std_logic_vector(to_unsigned( 247, 8)),
16 => std_logic_vector(to_unsigned( 97, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 272 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 58, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 89, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 176, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 114, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 51, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 198, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 70, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 273 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 136, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 34, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 36, 8)),
11 => std_logic_vector(to_unsigned( 236, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 34, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001011
elsif count = 274 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 237, 8)),
5 => std_logic_vector(to_unsigned( 43, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 64, 8)),
8 => std_logic_vector(to_unsigned( 244, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 95, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 138, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 275 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 153, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 51, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 55, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 49, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 78, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 276 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 102, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 177, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 177, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 244, 8)),
12 => std_logic_vector(to_unsigned( 196, 8)),
13 => std_logic_vector(to_unsigned( 228, 8)),
14 => std_logic_vector(to_unsigned( 214, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 197, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 277 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 71, 8)),
3 => std_logic_vector(to_unsigned( 181, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 35, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 57, 8)),
9 => std_logic_vector(to_unsigned( 21, 8)),
10 => std_logic_vector(to_unsigned( 242, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 243, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 68, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 278 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 143, 8)),
2 => std_logic_vector(to_unsigned( 225, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 198, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 131, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 84, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 182, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 279 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 244, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 235, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 31, 8)),
11 => std_logic_vector(to_unsigned( 163, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 67, 8)),
15 => std_logic_vector(to_unsigned( 9, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 280 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 33, 8)),
4 => std_logic_vector(to_unsigned( 239, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 28, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 34, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 77, 8)),
13 => std_logic_vector(to_unsigned( 185, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 57, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 281 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 192, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 216, 8)),
9 => std_logic_vector(to_unsigned( 138, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 110, 8)),
13 => std_logic_vector(to_unsigned( 94, 8)),
14 => std_logic_vector(to_unsigned( 63, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 282 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 24, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 61, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 76, 8)),
11 => std_logic_vector(to_unsigned( 34, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 45, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 71, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 283 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 251, 8)),
5 => std_logic_vector(to_unsigned( 243, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 244, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 284 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 162, 8)),
2 => std_logic_vector(to_unsigned( 22, 8)),
3 => std_logic_vector(to_unsigned( 39, 8)),
4 => std_logic_vector(to_unsigned( 232, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 188, 8)),
8 => std_logic_vector(to_unsigned( 251, 8)),
9 => std_logic_vector(to_unsigned( 141, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 188, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 285 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 130, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 26, 8)),
16 => std_logic_vector(to_unsigned( 63, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 286 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 40, 8)),
3 => std_logic_vector(to_unsigned( 15, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 110, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 2, 8)),
8 => std_logic_vector(to_unsigned( 83, 8)),
9 => std_logic_vector(to_unsigned( 229, 8)),
10 => std_logic_vector(to_unsigned( 177, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 243, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 18, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 287 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 121, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 83, 8)),
7 => std_logic_vector(to_unsigned( 101, 8)),
8 => std_logic_vector(to_unsigned( 182, 8)),
9 => std_logic_vector(to_unsigned( 243, 8)),
10 => std_logic_vector(to_unsigned( 36, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 172, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 29, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 288 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 150, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 63, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 133, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 214, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 157, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 289 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 3, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 95, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 190, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 290 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 216, 8)),
3 => std_logic_vector(to_unsigned( 120, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 223, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 76, 8)),
10 => std_logic_vector(to_unsigned( 210, 8)),
11 => std_logic_vector(to_unsigned( 28, 8)),
12 => std_logic_vector(to_unsigned( 250, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 202, 8)),
15 => std_logic_vector(to_unsigned( 39, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 291 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 156, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 104, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 247, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 292 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 176, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 219, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 208, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 293 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 212, 8)),
2 => std_logic_vector(to_unsigned( 115, 8)),
3 => std_logic_vector(to_unsigned( 196, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 74, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 224, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 159, 8)),
12 => std_logic_vector(to_unsigned( 20, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 228, 8)),
15 => std_logic_vector(to_unsigned( 63, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 294 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 198, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 222, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 132, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 250, 8)),
12 => std_logic_vector(to_unsigned( 206, 8)),
13 => std_logic_vector(to_unsigned( 195, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 48, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 295 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 236, 8)),
2 => std_logic_vector(to_unsigned( 59, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 84, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 10, 8)),
12 => std_logic_vector(to_unsigned( 43, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 237, 8)),
16 => std_logic_vector(to_unsigned( 162, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 296 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 55, 8)),
5 => std_logic_vector(to_unsigned( 101, 8)),
6 => std_logic_vector(to_unsigned( 45, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 36, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 193, 8)),
12 => std_logic_vector(to_unsigned( 185, 8)),
13 => std_logic_vector(to_unsigned( 176, 8)),
14 => std_logic_vector(to_unsigned( 41, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 49, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 62, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 297 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 221, 8)),
2 => std_logic_vector(to_unsigned( 94, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 28, 8)),
5 => std_logic_vector(to_unsigned( 205, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 207, 8)),
9 => std_logic_vector(to_unsigned( 28, 8)),
10 => std_logic_vector(to_unsigned( 180, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 74, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 83, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 298 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 240, 8)),
4 => std_logic_vector(to_unsigned( 55, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 250, 8)),
12 => std_logic_vector(to_unsigned( 5, 8)),
13 => std_logic_vector(to_unsigned( 232, 8)),
14 => std_logic_vector(to_unsigned( 233, 8)),
15 => std_logic_vector(to_unsigned( 180, 8)),
16 => std_logic_vector(to_unsigned( 64, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 299 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 223, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 222, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 179, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 155, 8)),
14 => std_logic_vector(to_unsigned( 244, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 207, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 300 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 232, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 249, 8)),
4 => std_logic_vector(to_unsigned( 102, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 191, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 237, 8)),
13 => std_logic_vector(to_unsigned( 33, 8)),
14 => std_logic_vector(to_unsigned( 146, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 301 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 30, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 90, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 197, 8)),
6 => std_logic_vector(to_unsigned( 202, 8)),
7 => std_logic_vector(to_unsigned( 91, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 100, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 241, 8)),
13 => std_logic_vector(to_unsigned( 33, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 302 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 208, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 150, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 1, 8)),
6 => std_logic_vector(to_unsigned( 182, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 112, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 31, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 303 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 0, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 210, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 228, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 187, 8)),
13 => std_logic_vector(to_unsigned( 176, 8)),
14 => std_logic_vector(to_unsigned( 57, 8)),
15 => std_logic_vector(to_unsigned( 2, 8)),
16 => std_logic_vector(to_unsigned( 241, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 304 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 195, 8)),
4 => std_logic_vector(to_unsigned( 173, 8)),
5 => std_logic_vector(to_unsigned( 5, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 96, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 173, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 305 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 185, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 107, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 190, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 32, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 213, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 306 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 65, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 166, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 119, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 50, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 307 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 42, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 158, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 56, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 84, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 191, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 308 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 29, 8)),
2 => std_logic_vector(to_unsigned( 227, 8)),
3 => std_logic_vector(to_unsigned( 214, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 137, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 196, 8)),
13 => std_logic_vector(to_unsigned( 176, 8)),
14 => std_logic_vector(to_unsigned( 15, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 309 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 181, 8)),
5 => std_logic_vector(to_unsigned( 38, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 100, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 96, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 234, 8)),
16 => std_logic_vector(to_unsigned( 7, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 310 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 226, 8)),
2 => std_logic_vector(to_unsigned( 23, 8)),
3 => std_logic_vector(to_unsigned( 31, 8)),
4 => std_logic_vector(to_unsigned( 245, 8)),
5 => std_logic_vector(to_unsigned( 240, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 204, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 99, 8)),
10 => std_logic_vector(to_unsigned( 239, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 175, 8)),
14 => std_logic_vector(to_unsigned( 52, 8)),
15 => std_logic_vector(to_unsigned( 241, 8)),
16 => std_logic_vector(to_unsigned( 54, 8)),
17 => std_logic_vector(to_unsigned( 209, 8)),
18 => std_logic_vector(to_unsigned( 46, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 311 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 163, 8)),
2 => std_logic_vector(to_unsigned( 208, 8)),
3 => std_logic_vector(to_unsigned( 101, 8)),
4 => std_logic_vector(to_unsigned( 30, 8)),
5 => std_logic_vector(to_unsigned( 161, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 181, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 206, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 18, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 312 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 55, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 50, 8)),
4 => std_logic_vector(to_unsigned( 37, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 233, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 196, 8)),
13 => std_logic_vector(to_unsigned( 241, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 44, 8)),
16 => std_logic_vector(to_unsigned( 249, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111100
elsif count = 313 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 89, 8)),
8 => std_logic_vector(to_unsigned( 132, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 27, 8)),
12 => std_logic_vector(to_unsigned( 16, 8)),
13 => std_logic_vector(to_unsigned( 138, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 314 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 213, 8)),
7 => std_logic_vector(to_unsigned( 180, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 137, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 135, 8)),
15 => std_logic_vector(to_unsigned( 6, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 315 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 229, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 171, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 212, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 4, 8)),
14 => std_logic_vector(to_unsigned( 238, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 316 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 185, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 30, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 95, 8)),
7 => std_logic_vector(to_unsigned( 174, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 9, 8)),
16 => std_logic_vector(to_unsigned( 20, 8)),
17 => std_logic_vector(to_unsigned( 196, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 317 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 111, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 212, 8)),
6 => std_logic_vector(to_unsigned( 172, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 224, 8)),
11 => std_logic_vector(to_unsigned( 228, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 250, 8)),
14 => std_logic_vector(to_unsigned( 79, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 318 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 75, 8)),
4 => std_logic_vector(to_unsigned( 79, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 204, 8)),
8 => std_logic_vector(to_unsigned( 250, 8)),
9 => std_logic_vector(to_unsigned( 80, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 235, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 214, 8)),
16 => std_logic_vector(to_unsigned( 11, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010111
elsif count = 319 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 17, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 19, 8)),
7 => std_logic_vector(to_unsigned( 71, 8)),
8 => std_logic_vector(to_unsigned( 221, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 215, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 232, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011000
elsif count = 320 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 61, 8)),
2 => std_logic_vector(to_unsigned( 246, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 207, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 62, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 44, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110110
elsif count = 321 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 33, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 239, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 61, 8)),
6 => std_logic_vector(to_unsigned( 88, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 86, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 191, 8)),
12 => std_logic_vector(to_unsigned( 2, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 126, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 322 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 10, 8)),
2 => std_logic_vector(to_unsigned( 32, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 54, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 183, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 130, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 177, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 226, 8)),
13 => std_logic_vector(to_unsigned( 36, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 323 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 194, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 37, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 8, 8)),
8 => std_logic_vector(to_unsigned( 165, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 155, 8)),
14 => std_logic_vector(to_unsigned( 220, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 74, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010011
elsif count = 324 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 159, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 243, 8)),
12 => std_logic_vector(to_unsigned( 216, 8)),
13 => std_logic_vector(to_unsigned( 201, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 149, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 325 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 27, 8)),
4 => std_logic_vector(to_unsigned( 240, 8)),
5 => std_logic_vector(to_unsigned( 232, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 21, 8)),
8 => std_logic_vector(to_unsigned( 89, 8)),
9 => std_logic_vector(to_unsigned( 41, 8)),
10 => std_logic_vector(to_unsigned( 156, 8)),
11 => std_logic_vector(to_unsigned( 72, 8)),
12 => std_logic_vector(to_unsigned( 187, 8)),
13 => std_logic_vector(to_unsigned( 79, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 29, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 326 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 75, 8)),
3 => std_logic_vector(to_unsigned( 224, 8)),
4 => std_logic_vector(to_unsigned( 254, 8)),
5 => std_logic_vector(to_unsigned( 190, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 173, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 21, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 102, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 327 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 77, 8)),
2 => std_logic_vector(to_unsigned( 164, 8)),
3 => std_logic_vector(to_unsigned( 9, 8)),
4 => std_logic_vector(to_unsigned( 18, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 192, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 183, 8)),
12 => std_logic_vector(to_unsigned( 198, 8)),
13 => std_logic_vector(to_unsigned( 212, 8)),
14 => std_logic_vector(to_unsigned( 130, 8)),
15 => std_logic_vector(to_unsigned( 239, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 328 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 18, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 25, 8)),
7 => std_logic_vector(to_unsigned( 98, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 95, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 42, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 78, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 329 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 59, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 130, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 210, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 73, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 330 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 229, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 171, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 23, 8)),
11 => std_logic_vector(to_unsigned( 208, 8)),
12 => std_logic_vector(to_unsigned( 20, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 50, 8)),
15 => std_logic_vector(to_unsigned( 90, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 51, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000110
elsif count = 331 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 42, 8)),
3 => std_logic_vector(to_unsigned( 41, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 43, 8)),
8 => std_logic_vector(to_unsigned( 77, 8)),
9 => std_logic_vector(to_unsigned( 41, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 134, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 332 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 35, 8)),
8 => std_logic_vector(to_unsigned( 214, 8)),
9 => std_logic_vector(to_unsigned( 255, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 191, 8)),
12 => std_logic_vector(to_unsigned( 145, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 238, 8)),
16 => std_logic_vector(to_unsigned( 162, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 333 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 198, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 183, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 230, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 187, 8)),
16 => std_logic_vector(to_unsigned( 236, 8)),
17 => std_logic_vector(to_unsigned( 196, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 334 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 219, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 218, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 193, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 224, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 335 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 210, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 187, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 229, 8)),
7 => std_logic_vector(to_unsigned( 15, 8)),
8 => std_logic_vector(to_unsigned( 218, 8)),
9 => std_logic_vector(to_unsigned( 233, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 10, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 185, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 336 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 17, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 72, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 33, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 133, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 337 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 78, 8)),
8 => std_logic_vector(to_unsigned( 213, 8)),
9 => std_logic_vector(to_unsigned( 230, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 151, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 86, 8)),
16 => std_logic_vector(to_unsigned( 207, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 338 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 136, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 9, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 35, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 36, 8)),
9 => std_logic_vector(to_unsigned( 53, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 255, 8)),
13 => std_logic_vector(to_unsigned( 37, 8)),
14 => std_logic_vector(to_unsigned( 50, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 70, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 339 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 182, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 202, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 229, 8)),
8 => std_logic_vector(to_unsigned( 131, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 203, 8)),
11 => std_logic_vector(to_unsigned( 136, 8)),
12 => std_logic_vector(to_unsigned( 226, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 340 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 11, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 195, 8)),
5 => std_logic_vector(to_unsigned( 163, 8)),
6 => std_logic_vector(to_unsigned( 238, 8)),
7 => std_logic_vector(to_unsigned( 251, 8)),
8 => std_logic_vector(to_unsigned( 12, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 239, 8)),
11 => std_logic_vector(to_unsigned( 213, 8)),
12 => std_logic_vector(to_unsigned( 203, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 246, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 341 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 221, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 208, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 246, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 246, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 228, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 0, 8)),
17 => std_logic_vector(to_unsigned( 218, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 342 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 37, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 20, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 12, 8)),
11 => std_logic_vector(to_unsigned( 43, 8)),
12 => std_logic_vector(to_unsigned( 46, 8)),
13 => std_logic_vector(to_unsigned( 28, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 343 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 151, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 43, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 16, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 165, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 200, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 56, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 344 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 230, 8)),
4 => std_logic_vector(to_unsigned( 63, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 71, 8)),
7 => std_logic_vector(to_unsigned( 24, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 21, 8)),
10 => std_logic_vector(to_unsigned( 245, 8)),
11 => std_logic_vector(to_unsigned( 234, 8)),
12 => std_logic_vector(to_unsigned( 57, 8)),
13 => std_logic_vector(to_unsigned( 185, 8)),
14 => std_logic_vector(to_unsigned( 10, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 24, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 58, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 345 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 32, 8)),
7 => std_logic_vector(to_unsigned( 48, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 157, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 116, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 346 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 148, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 217, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 199, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 13, 8)),
10 => std_logic_vector(to_unsigned( 251, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 34, 8)),
14 => std_logic_vector(to_unsigned( 37, 8)),
15 => std_logic_vector(to_unsigned( 187, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100110
elsif count = 347 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 62, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 187, 8)),
5 => std_logic_vector(to_unsigned( 29, 8)),
6 => std_logic_vector(to_unsigned( 33, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 118, 8)),
10 => std_logic_vector(to_unsigned( 245, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 244, 8)),
13 => std_logic_vector(to_unsigned( 7, 8)),
14 => std_logic_vector(to_unsigned( 23, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 254, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111010
elsif count = 348 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 95, 8)),
2 => std_logic_vector(to_unsigned( 21, 8)),
3 => std_logic_vector(to_unsigned( 233, 8)),
4 => std_logic_vector(to_unsigned( 9, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 140, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 78, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 349 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 68, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 7, 8)),
7 => std_logic_vector(to_unsigned( 173, 8)),
8 => std_logic_vector(to_unsigned( 216, 8)),
9 => std_logic_vector(to_unsigned( 200, 8)),
10 => std_logic_vector(to_unsigned( 221, 8)),
11 => std_logic_vector(to_unsigned( 159, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 95, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 350 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 175, 8)),
3 => std_logic_vector(to_unsigned( 169, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 241, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 217, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 20, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 227, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 86, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 351 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 2, 8)),
5 => std_logic_vector(to_unsigned( 189, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 79, 8)),
11 => std_logic_vector(to_unsigned( 188, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 190, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 352 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 117, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 193, 8)),
7 => std_logic_vector(to_unsigned( 233, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 248, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 138, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 45, 8)),
16 => std_logic_vector(to_unsigned( 45, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 353 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 162, 8)),
2 => std_logic_vector(to_unsigned( 91, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 73, 8)),
5 => std_logic_vector(to_unsigned( 41, 8)),
6 => std_logic_vector(to_unsigned( 159, 8)),
7 => std_logic_vector(to_unsigned( 57, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 138, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 154, 8)),
16 => std_logic_vector(to_unsigned( 153, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 354 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 136, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 198, 8)),
6 => std_logic_vector(to_unsigned( 212, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 184, 8)),
10 => std_logic_vector(to_unsigned( 64, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 103, 8)),
16 => std_logic_vector(to_unsigned( 80, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 355 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 63, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 243, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 90, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 126, 8)),
15 => std_logic_vector(to_unsigned( 74, 8)),
16 => std_logic_vector(to_unsigned( 5, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 356 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 48, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 53, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 67, 8)),
8 => std_logic_vector(to_unsigned( 51, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 86, 8)),
13 => std_logic_vector(to_unsigned( 237, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 139, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 357 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 178, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 51, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 180, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 126, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 206, 8)),
12 => std_logic_vector(to_unsigned( 173, 8)),
13 => std_logic_vector(to_unsigned( 213, 8)),
14 => std_logic_vector(to_unsigned( 179, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 358 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 158, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 16, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 33, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 26, 8)),
15 => std_logic_vector(to_unsigned( 55, 8)),
16 => std_logic_vector(to_unsigned( 77, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 359 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 208, 8)),
2 => std_logic_vector(to_unsigned( 57, 8)),
3 => std_logic_vector(to_unsigned( 237, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 7, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 245, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 216, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 360 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 235, 8)),
2 => std_logic_vector(to_unsigned( 0, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 207, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 228, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 230, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 211, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 211, 8)),
17 => std_logic_vector(to_unsigned( 51, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 361 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 16, 8)),
2 => std_logic_vector(to_unsigned( 84, 8)),
3 => std_logic_vector(to_unsigned( 178, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 183, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 103, 8)),
8 => std_logic_vector(to_unsigned( 59, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 139, 8)),
11 => std_logic_vector(to_unsigned( 218, 8)),
12 => std_logic_vector(to_unsigned( 168, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 362 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 182, 8)),
6 => std_logic_vector(to_unsigned( 172, 8)),
7 => std_logic_vector(to_unsigned( 1, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 215, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 213, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 247, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 205, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110011
elsif count = 363 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 192, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 249, 8)),
7 => std_logic_vector(to_unsigned( 71, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 13, 8)),
10 => std_logic_vector(to_unsigned( 221, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 230, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 230, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 123, 8)),
18 => std_logic_vector(to_unsigned( 193, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 364 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 211, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 45, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 44, 8)),
13 => std_logic_vector(to_unsigned( 180, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 6, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 365 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 5, 8)),
2 => std_logic_vector(to_unsigned( 197, 8)),
3 => std_logic_vector(to_unsigned( 150, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 123, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 215, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 31, 8)),
16 => std_logic_vector(to_unsigned( 14, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 366 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 55, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 70, 8)),
4 => std_logic_vector(to_unsigned( 185, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 136, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 181, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 9, 8)),
13 => std_logic_vector(to_unsigned( 156, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 132, 8)),
16 => std_logic_vector(to_unsigned( 145, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 367 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 34, 8)),
4 => std_logic_vector(to_unsigned( 242, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 134, 8)),
7 => std_logic_vector(to_unsigned( 249, 8)),
8 => std_logic_vector(to_unsigned( 22, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 368 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 60, 8)),
2 => std_logic_vector(to_unsigned( 155, 8)),
3 => std_logic_vector(to_unsigned( 159, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 189, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 212, 8)),
8 => std_logic_vector(to_unsigned( 164, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 213, 8)),
12 => std_logic_vector(to_unsigned( 163, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 369 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 63, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 242, 8)),
6 => std_logic_vector(to_unsigned( 11, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 89, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 121, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 370 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 18, 8)),
2 => std_logic_vector(to_unsigned( 185, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 59, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 251, 8)),
9 => std_logic_vector(to_unsigned( 24, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 237, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 193, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001101
elsif count = 371 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 235, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 137, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 153, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 234, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 217, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 207, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 372 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 232, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 62, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 4, 8)),
8 => std_logic_vector(to_unsigned( 95, 8)),
9 => std_logic_vector(to_unsigned( 204, 8)),
10 => std_logic_vector(to_unsigned( 144, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 173, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 192, 8)),
16 => std_logic_vector(to_unsigned( 156, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 373 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 4, 8)),
2 => std_logic_vector(to_unsigned( 175, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 24, 8)),
8 => std_logic_vector(to_unsigned( 155, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 177, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 140, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 12, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 374 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 14, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 144, 8)),
9 => std_logic_vector(to_unsigned( 23, 8)),
10 => std_logic_vector(to_unsigned( 56, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 237, 8)),
13 => std_logic_vector(to_unsigned( 188, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 375 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 143, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 112, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 145, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 376 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 22, 8)),
3 => std_logic_vector(to_unsigned( 20, 8)),
4 => std_logic_vector(to_unsigned( 59, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 219, 8)),
10 => std_logic_vector(to_unsigned( 16, 8)),
11 => std_logic_vector(to_unsigned( 56, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 213, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 210, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 377 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 136, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 238, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 94, 8)),
7 => std_logic_vector(to_unsigned( 236, 8)),
8 => std_logic_vector(to_unsigned( 74, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 61, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 188, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 378 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 177, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 43, 8)),
5 => std_logic_vector(to_unsigned( 17, 8)),
6 => std_logic_vector(to_unsigned( 34, 8)),
7 => std_logic_vector(to_unsigned( 22, 8)),
8 => std_logic_vector(to_unsigned( 137, 8)),
9 => std_logic_vector(to_unsigned( 174, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 100, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 53, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 24, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 379 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 0, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 11, 8)),
4 => std_logic_vector(to_unsigned( 62, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 189, 8)),
9 => std_logic_vector(to_unsigned( 238, 8)),
10 => std_logic_vector(to_unsigned( 3, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 232, 8)),
13 => std_logic_vector(to_unsigned( 154, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 380 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 55, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 151, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 381 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 80, 8)),
2 => std_logic_vector(to_unsigned( 39, 8)),
3 => std_logic_vector(to_unsigned( 174, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 12, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 69, 8)),
9 => std_logic_vector(to_unsigned( 30, 8)),
10 => std_logic_vector(to_unsigned( 59, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 17, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 17, 8)),
15 => std_logic_vector(to_unsigned( 227, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 53, 8)),
18 => std_logic_vector(to_unsigned( 47, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 382 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 128, 8)),
2 => std_logic_vector(to_unsigned( 54, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 47, 8)),
5 => std_logic_vector(to_unsigned( 209, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 23, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 64, 8)),
11 => std_logic_vector(to_unsigned( 142, 8)),
12 => std_logic_vector(to_unsigned( 88, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 31, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 26, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 53, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 383 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 254, 8)),
2 => std_logic_vector(to_unsigned( 206, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 13, 8)),
8 => std_logic_vector(to_unsigned( 37, 8)),
9 => std_logic_vector(to_unsigned( 234, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 229, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 73, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 58, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 384 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 24, 8)),
2 => std_logic_vector(to_unsigned( 157, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 177, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 236, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 201, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 234, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 385 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 238, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 115, 8)),
7 => std_logic_vector(to_unsigned( 209, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 76, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 46, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 152, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110110
elsif count = 386 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 75, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 184, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 37, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 21, 8)),
14 => std_logic_vector(to_unsigned( 165, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 387 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 163, 8)),
2 => std_logic_vector(to_unsigned( 33, 8)),
3 => std_logic_vector(to_unsigned( 165, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 25, 8)),
6 => std_logic_vector(to_unsigned( 218, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 52, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 105, 8)),
14 => std_logic_vector(to_unsigned( 235, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 56, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 388 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 143, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 254, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 244, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 159, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 136, 8)),
14 => std_logic_vector(to_unsigned( 140, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 389 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 130, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 14, 8)),
5 => std_logic_vector(to_unsigned( 216, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 20, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 207, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 60, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 390 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 59, 8)),
2 => std_logic_vector(to_unsigned( 90, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 89, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 27, 8)),
8 => std_logic_vector(to_unsigned( 58, 8)),
9 => std_logic_vector(to_unsigned( 29, 8)),
10 => std_logic_vector(to_unsigned( 54, 8)),
11 => std_logic_vector(to_unsigned( 0, 8)),
12 => std_logic_vector(to_unsigned( 186, 8)),
13 => std_logic_vector(to_unsigned( 156, 8)),
14 => std_logic_vector(to_unsigned( 62, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 59, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 391 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 25, 8)),
2 => std_logic_vector(to_unsigned( 202, 8)),
3 => std_logic_vector(to_unsigned( 166, 8)),
4 => std_logic_vector(to_unsigned( 79, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 152, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 90, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 128, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 392 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 231, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 46, 8)),
6 => std_logic_vector(to_unsigned( 137, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 110, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 78, 8)),
12 => std_logic_vector(to_unsigned( 105, 8)),
13 => std_logic_vector(to_unsigned( 185, 8)),
14 => std_logic_vector(to_unsigned( 16, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 393 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 160, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 82, 8)),
6 => std_logic_vector(to_unsigned( 154, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 204, 8)),
9 => std_logic_vector(to_unsigned( 0, 8)),
10 => std_logic_vector(to_unsigned( 136, 8)),
11 => std_logic_vector(to_unsigned( 19, 8)),
12 => std_logic_vector(to_unsigned( 255, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 194, 8)),
15 => std_logic_vector(to_unsigned( 113, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 394 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 59, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 37, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 113, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 181, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 137, 8)),
11 => std_logic_vector(to_unsigned( 17, 8)),
12 => std_logic_vector(to_unsigned( 210, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 61, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 395 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 247, 8)),
2 => std_logic_vector(to_unsigned( 238, 8)),
3 => std_logic_vector(to_unsigned( 159, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 95, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 103, 8)),
10 => std_logic_vector(to_unsigned( 166, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 192, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 396 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 147, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 247, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 138, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 151, 8)),
14 => std_logic_vector(to_unsigned( 158, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 397 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 149, 8)),
4 => std_logic_vector(to_unsigned( 170, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 28, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 63, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 123, 8)),
16 => std_logic_vector(to_unsigned( 203, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 398 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 186, 8)),
4 => std_logic_vector(to_unsigned( 91, 8)),
5 => std_logic_vector(to_unsigned( 148, 8)),
6 => std_logic_vector(to_unsigned( 11, 8)),
7 => std_logic_vector(to_unsigned( 2, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 14, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 139, 8)),
18 => std_logic_vector(to_unsigned( 70, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 399 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 141, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 230, 8)),
5 => std_logic_vector(to_unsigned( 180, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 66, 8)),
10 => std_logic_vector(to_unsigned( 206, 8)),
11 => std_logic_vector(to_unsigned( 211, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 194, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 400 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 186, 8)),
4 => std_logic_vector(to_unsigned( 80, 8)),
5 => std_logic_vector(to_unsigned( 180, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 85, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 90, 8)),
13 => std_logic_vector(to_unsigned( 141, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 51, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 61, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 401 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 27, 8)),
2 => std_logic_vector(to_unsigned( 14, 8)),
3 => std_logic_vector(to_unsigned( 90, 8)),
4 => std_logic_vector(to_unsigned( 207, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 86, 8)),
10 => std_logic_vector(to_unsigned( 200, 8)),
11 => std_logic_vector(to_unsigned( 188, 8)),
12 => std_logic_vector(to_unsigned( 188, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 86, 8)),
16 => std_logic_vector(to_unsigned( 253, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 402 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 220, 8)),
3 => std_logic_vector(to_unsigned( 26, 8)),
4 => std_logic_vector(to_unsigned( 244, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 14, 8)),
11 => std_logic_vector(to_unsigned( 92, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 135, 8)),
14 => std_logic_vector(to_unsigned( 231, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 403 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 22, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 14, 8)),
4 => std_logic_vector(to_unsigned( 20, 8)),
5 => std_logic_vector(to_unsigned( 44, 8)),
6 => std_logic_vector(to_unsigned( 45, 8)),
7 => std_logic_vector(to_unsigned( 207, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 11, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 36, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 18, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100100
elsif count = 404 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 34, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 50, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 58, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 108, 8)),
11 => std_logic_vector(to_unsigned( 200, 8)),
12 => std_logic_vector(to_unsigned( 233, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010101
elsif count = 405 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 99, 8)),
2 => std_logic_vector(to_unsigned( 243, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 60, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 13, 8)),
10 => std_logic_vector(to_unsigned( 122, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 249, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 68, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 406 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 69, 8)),
2 => std_logic_vector(to_unsigned( 223, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 22, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 188, 8)),
10 => std_logic_vector(to_unsigned( 136, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 48, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 191, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 407 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 141, 8)),
2 => std_logic_vector(to_unsigned( 88, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 79, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 89, 8)),
9 => std_logic_vector(to_unsigned( 176, 8)),
10 => std_logic_vector(to_unsigned( 254, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 227, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 408 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 244, 8)),
4 => std_logic_vector(to_unsigned( 185, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 140, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 47, 8)),
15 => std_logic_vector(to_unsigned( 247, 8)),
16 => std_logic_vector(to_unsigned( 217, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 58, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 409 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 212, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 227, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 235, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 36, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 174, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 410 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 120, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 17, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 166, 8)),
16 => std_logic_vector(to_unsigned( 55, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 411 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 160, 8)),
3 => std_logic_vector(to_unsigned( 91, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 31, 8)),
6 => std_logic_vector(to_unsigned( 251, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 177, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 412 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 244, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 209, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 237, 8)),
10 => std_logic_vector(to_unsigned( 182, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 227, 8)),
13 => std_logic_vector(to_unsigned( 39, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 56, 8)),
16 => std_logic_vector(to_unsigned( 202, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 413 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 111, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 230, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 52, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 42, 8)),
14 => std_logic_vector(to_unsigned( 57, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 98, 8)),
17 => std_logic_vector(to_unsigned( 59, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 414 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 61, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 200, 8)),
7 => std_logic_vector(to_unsigned( 154, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 159, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 48, 8)),
16 => std_logic_vector(to_unsigned( 36, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 415 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 185, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 171, 8)),
4 => std_logic_vector(to_unsigned( 22, 8)),
5 => std_logic_vector(to_unsigned( 207, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 17, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 16, 8)),
11 => std_logic_vector(to_unsigned( 249, 8)),
12 => std_logic_vector(to_unsigned( 185, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 2, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 39, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 416 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 52, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 18, 8)),
6 => std_logic_vector(to_unsigned( 62, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 130, 8)),
9 => std_logic_vector(to_unsigned( 57, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 41, 8)),
13 => std_logic_vector(to_unsigned( 150, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 417 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 187, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 188, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 103, 8)),
7 => std_logic_vector(to_unsigned( 39, 8)),
8 => std_logic_vector(to_unsigned( 166, 8)),
9 => std_logic_vector(to_unsigned( 200, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 150, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 418 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 81, 8)),
2 => std_logic_vector(to_unsigned( 221, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 237, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 50, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 217, 8)),
15 => std_logic_vector(to_unsigned( 251, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 419 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 12, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 238, 8)),
5 => std_logic_vector(to_unsigned( 51, 8)),
6 => std_logic_vector(to_unsigned( 60, 8)),
7 => std_logic_vector(to_unsigned( 172, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 242, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 203, 8)),
15 => std_logic_vector(to_unsigned( 237, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 47, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110011
elsif count = 420 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 170, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 214, 8)),
9 => std_logic_vector(to_unsigned( 33, 8)),
10 => std_logic_vector(to_unsigned( 56, 8)),
11 => std_logic_vector(to_unsigned( 132, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 421 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 177, 8)),
3 => std_logic_vector(to_unsigned( 56, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 17, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 136, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 187, 8)),
13 => std_logic_vector(to_unsigned( 80, 8)),
14 => std_logic_vector(to_unsigned( 1, 8)),
15 => std_logic_vector(to_unsigned( 18, 8)),
16 => std_logic_vector(to_unsigned( 183, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 181, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 422 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 212, 8)),
2 => std_logic_vector(to_unsigned( 190, 8)),
3 => std_logic_vector(to_unsigned( 230, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 180, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 185, 8)),
9 => std_logic_vector(to_unsigned( 134, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 35, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 177, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 423 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 54, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 151, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 244, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 213, 8)),
14 => std_logic_vector(to_unsigned( 135, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 73, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 424 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 216, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 52, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 31, 8)),
10 => std_logic_vector(to_unsigned( 189, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 72, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 425 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 78, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 132, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 214, 8)),
10 => std_logic_vector(to_unsigned( 68, 8)),
11 => std_logic_vector(to_unsigned( 124, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 181, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 241, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 426 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 166, 8)),
2 => std_logic_vector(to_unsigned( 84, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 209, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 236, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 186, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 203, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 427 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 82, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 32, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 194, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 92, 8)),
11 => std_logic_vector(to_unsigned( 60, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 135, 8)),
14 => std_logic_vector(to_unsigned( 182, 8)),
15 => std_logic_vector(to_unsigned( 99, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 128, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 428 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 12, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 63, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 156, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 140, 8)),
11 => std_logic_vector(to_unsigned( 7, 8)),
12 => std_logic_vector(to_unsigned( 230, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 163, 8)),
15 => std_logic_vector(to_unsigned( 19, 8)),
16 => std_logic_vector(to_unsigned( 156, 8)),
17 => std_logic_vector(to_unsigned( 51, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 429 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 204, 8)),
2 => std_logic_vector(to_unsigned( 8, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 148, 8)),
6 => std_logic_vector(to_unsigned( 192, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 222, 8)),
11 => std_logic_vector(to_unsigned( 72, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 226, 8)),
14 => std_logic_vector(to_unsigned( 37, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 185, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 430 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 55, 8)),
2 => std_logic_vector(to_unsigned( 246, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 159, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 210, 8)),
12 => std_logic_vector(to_unsigned( 203, 8)),
13 => std_logic_vector(to_unsigned( 151, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 253, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 431 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 254, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 17, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 104, 8)),
9 => std_logic_vector(to_unsigned( 19, 8)),
10 => std_logic_vector(to_unsigned( 3, 8)),
11 => std_logic_vector(to_unsigned( 65, 8)),
12 => std_logic_vector(to_unsigned( 109, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 75, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 78, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101010
elsif count = 432 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 79, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 224, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 95, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 433 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 223, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 209, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 213, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 230, 8)),
12 => std_logic_vector(to_unsigned( 208, 8)),
13 => std_logic_vector(to_unsigned( 150, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 231, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 434 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 41, 8)),
2 => std_logic_vector(to_unsigned( 255, 8)),
3 => std_logic_vector(to_unsigned( 252, 8)),
4 => std_logic_vector(to_unsigned( 91, 8)),
5 => std_logic_vector(to_unsigned( 14, 8)),
6 => std_logic_vector(to_unsigned( 12, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 151, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 60, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 97, 8)),
17 => std_logic_vector(to_unsigned( 52, 8)),
18 => std_logic_vector(to_unsigned( 106, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 435 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 63, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 209, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 250, 8)),
11 => std_logic_vector(to_unsigned( 206, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 37, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 60, 8)),
17 => std_logic_vector(to_unsigned( 139, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 436 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 196, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 44, 8)),
6 => std_logic_vector(to_unsigned( 30, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 80, 8)),
10 => std_logic_vector(to_unsigned( 12, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 51, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 63, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 437 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 249, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 220, 8)),
7 => std_logic_vector(to_unsigned( 56, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 222, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 438 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 54, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 78, 8)),
5 => std_logic_vector(to_unsigned( 26, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 63, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 232, 8)),
10 => std_logic_vector(to_unsigned( 223, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 66, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 51, 8)),
15 => std_logic_vector(to_unsigned( 32, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 56, 8)),
18 => std_logic_vector(to_unsigned( 60, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 439 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 76, 8)),
2 => std_logic_vector(to_unsigned( 228, 8)),
3 => std_logic_vector(to_unsigned( 109, 8)),
4 => std_logic_vector(to_unsigned( 191, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 128, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 124, 8)),
11 => std_logic_vector(to_unsigned( 132, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 211, 8)),
15 => std_logic_vector(to_unsigned( 237, 8)),
16 => std_logic_vector(to_unsigned( 220, 8)),
17 => std_logic_vector(to_unsigned( 81, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 440 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 245, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 43, 8)),
7 => std_logic_vector(to_unsigned( 82, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 32, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 17, 8)),
15 => std_logic_vector(to_unsigned( 78, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 133, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 441 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 77, 8)),
2 => std_logic_vector(to_unsigned( 63, 8)),
3 => std_logic_vector(to_unsigned( 245, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 54, 8)),
8 => std_logic_vector(to_unsigned( 86, 8)),
9 => std_logic_vector(to_unsigned( 133, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 179, 8)),
13 => std_logic_vector(to_unsigned( 218, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 56, 8)),
16 => std_logic_vector(to_unsigned( 228, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 442 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 253, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 183, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 63, 8)),
10 => std_logic_vector(to_unsigned( 79, 8)),
11 => std_logic_vector(to_unsigned( 131, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 44, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 443 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 91, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 64, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 138, 8)),
11 => std_logic_vector(to_unsigned( 121, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 235, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 444 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 87, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 55, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 53, 8)),
6 => std_logic_vector(to_unsigned( 35, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 81, 8)),
9 => std_logic_vector(to_unsigned( 119, 8)),
10 => std_logic_vector(to_unsigned( 9, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 79, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 228, 8)),
16 => std_logic_vector(to_unsigned( 23, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 445 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 234, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 243, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 186, 8)),
9 => std_logic_vector(to_unsigned( 227, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 21, 8)),
13 => std_logic_vector(to_unsigned( 232, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 15, 8)),
17 => std_logic_vector(to_unsigned( 196, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 446 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 67, 8)),
3 => std_logic_vector(to_unsigned( 26, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 0, 8)),
6 => std_logic_vector(to_unsigned( 234, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 60, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 131, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 39, 8)),
13 => std_logic_vector(to_unsigned( 199, 8)),
14 => std_logic_vector(to_unsigned( 63, 8)),
15 => std_logic_vector(to_unsigned( 37, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 54, 8)),
18 => std_logic_vector(to_unsigned( 52, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 447 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 47, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 81, 8)),
4 => std_logic_vector(to_unsigned( 66, 8)),
5 => std_logic_vector(to_unsigned( 76, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 37, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 48, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 215, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 13, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 448 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 78, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 103, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 222, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 230, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 231, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 449 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 7, 8)),
6 => std_logic_vector(to_unsigned( 127, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 246, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 222, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 40, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 450 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 100, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 61, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 104, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 116, 8)),
11 => std_logic_vector(to_unsigned( 111, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 53, 8)),
14 => std_logic_vector(to_unsigned( 205, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 190, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 451 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 54, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 68, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 177, 8)),
10 => std_logic_vector(to_unsigned( 108, 8)),
11 => std_logic_vector(to_unsigned( 228, 8)),
12 => std_logic_vector(to_unsigned( 54, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 104, 8)),
16 => std_logic_vector(to_unsigned( 75, 8)),
17 => std_logic_vector(to_unsigned( 76, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 452 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 47, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 32, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 223, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 230, 8)),
12 => std_logic_vector(to_unsigned( 225, 8)),
13 => std_logic_vector(to_unsigned( 50, 8)),
14 => std_logic_vector(to_unsigned( 63, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 97, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 453 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 72, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 33, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 31, 8)),
11 => std_logic_vector(to_unsigned( 107, 8)),
12 => std_logic_vector(to_unsigned( 40, 8)),
13 => std_logic_vector(to_unsigned( 240, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 105, 8)),
17 => std_logic_vector(to_unsigned( 53, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 454 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 166, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 32, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 20, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 46, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 50, 8)),
13 => std_logic_vector(to_unsigned( 176, 8)),
14 => std_logic_vector(to_unsigned( 62, 8)),
15 => std_logic_vector(to_unsigned( 54, 8)),
16 => std_logic_vector(to_unsigned( 52, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 41, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 455 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 185, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 209, 8)),
7 => std_logic_vector(to_unsigned( 6, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 60, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 163, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 456 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 27, 8)),
2 => std_logic_vector(to_unsigned( 121, 8)),
3 => std_logic_vector(to_unsigned( 62, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 221, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 51, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 35, 8)),
13 => std_logic_vector(to_unsigned( 57, 8)),
14 => std_logic_vector(to_unsigned( 45, 8)),
15 => std_logic_vector(to_unsigned( 239, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 457 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 95, 8)),
5 => std_logic_vector(to_unsigned( 198, 8)),
6 => std_logic_vector(to_unsigned( 255, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 108, 8)),
11 => std_logic_vector(to_unsigned( 163, 8)),
12 => std_logic_vector(to_unsigned( 250, 8)),
13 => std_logic_vector(to_unsigned( 210, 8)),
14 => std_logic_vector(to_unsigned( 220, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 173, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 458 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 65, 8)),
2 => std_logic_vector(to_unsigned( 96, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 100, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 178, 8)),
11 => std_logic_vector(to_unsigned( 212, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 240, 8)),
14 => std_logic_vector(to_unsigned( 8, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 459 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 240, 8)),
3 => std_logic_vector(to_unsigned( 199, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 221, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 226, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 127, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 250, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 154, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 460 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 182, 8)),
3 => std_logic_vector(to_unsigned( 218, 8)),
4 => std_logic_vector(to_unsigned( 2, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 128, 8)),
8 => std_logic_vector(to_unsigned( 68, 8)),
9 => std_logic_vector(to_unsigned( 237, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 220, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 461 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 20, 8)),
8 => std_logic_vector(to_unsigned( 227, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 200, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 71, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 186, 8)),
15 => std_logic_vector(to_unsigned( 237, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 462 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 232, 8)),
5 => std_logic_vector(to_unsigned( 246, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 245, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 244, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 231, 8)),
15 => std_logic_vector(to_unsigned( 45, 8)),
16 => std_logic_vector(to_unsigned( 8, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 214, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 463 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 80, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 131, 8)),
9 => std_logic_vector(to_unsigned( 238, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 229, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 180, 8)),
14 => std_logic_vector(to_unsigned( 1, 8)),
15 => std_logic_vector(to_unsigned( 52, 8)),
16 => std_logic_vector(to_unsigned( 178, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101110
elsif count = 464 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 54, 8)),
2 => std_logic_vector(to_unsigned( 41, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 57, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 55, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 465 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 108, 8)),
4 => std_logic_vector(to_unsigned( 177, 8)),
5 => std_logic_vector(to_unsigned( 46, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 47, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 167, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 466 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 72, 8)),
5 => std_logic_vector(to_unsigned( 170, 8)),
6 => std_logic_vector(to_unsigned( 134, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 190, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 92, 8)),
16 => std_logic_vector(to_unsigned( 233, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 467 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 111, 8)),
2 => std_logic_vector(to_unsigned( 194, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 78, 8)),
6 => std_logic_vector(to_unsigned( 227, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 210, 8)),
9 => std_logic_vector(to_unsigned( 90, 8)),
10 => std_logic_vector(to_unsigned( 235, 8)),
11 => std_logic_vector(to_unsigned( 45, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 53, 8)),
14 => std_logic_vector(to_unsigned( 220, 8)),
15 => std_logic_vector(to_unsigned( 232, 8)),
16 => std_logic_vector(to_unsigned( 197, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 185, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 468 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 87, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 88, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 238, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 147, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 149, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101100
elsif count = 469 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 249, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 240, 8)),
7 => std_logic_vector(to_unsigned( 141, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 118, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 204, 8)),
12 => std_logic_vector(to_unsigned( 249, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 470 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 184, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 190, 8)),
10 => std_logic_vector(to_unsigned( 56, 8)),
11 => std_logic_vector(to_unsigned( 210, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 471 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 187, 8)),
3 => std_logic_vector(to_unsigned( 131, 8)),
4 => std_logic_vector(to_unsigned( 0, 8)),
5 => std_logic_vector(to_unsigned( 91, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 56, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 195, 8)),
11 => std_logic_vector(to_unsigned( 242, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 85, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 241, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001101
elsif count = 472 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 180, 8)),
2 => std_logic_vector(to_unsigned( 243, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 23, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 16, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 29, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 73, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011100
elsif count = 473 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 68, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 80, 8)),
5 => std_logic_vector(to_unsigned( 55, 8)),
6 => std_logic_vector(to_unsigned( 59, 8)),
7 => std_logic_vector(to_unsigned( 216, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 90, 8)),
10 => std_logic_vector(to_unsigned( 12, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 30, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 170, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 42, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 474 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 117, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 31, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 181, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 41, 8)),
13 => std_logic_vector(to_unsigned( 66, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 475 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 7, 8)),
3 => std_logic_vector(to_unsigned( 112, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 3, 8)),
7 => std_logic_vector(to_unsigned( 23, 8)),
8 => std_logic_vector(to_unsigned( 164, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 153, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 476 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 87, 8)),
2 => std_logic_vector(to_unsigned( 30, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 26, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 40, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 219, 8)),
15 => std_logic_vector(to_unsigned( 229, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 477 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 74, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 29, 8)),
4 => std_logic_vector(to_unsigned( 117, 8)),
5 => std_logic_vector(to_unsigned( 43, 8)),
6 => std_logic_vector(to_unsigned( 74, 8)),
7 => std_logic_vector(to_unsigned( 21, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 179, 8)),
11 => std_logic_vector(to_unsigned( 240, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 57, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 478 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 179, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 38, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 224, 8)),
8 => std_logic_vector(to_unsigned( 72, 8)),
9 => std_logic_vector(to_unsigned( 182, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 221, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 201, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 479 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 64, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 75, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 240, 8)),
12 => std_logic_vector(to_unsigned( 224, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 145, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 480 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 213, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 127, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 178, 8)),
11 => std_logic_vector(to_unsigned( 37, 8)),
12 => std_logic_vector(to_unsigned( 226, 8)),
13 => std_logic_vector(to_unsigned( 214, 8)),
14 => std_logic_vector(to_unsigned( 172, 8)),
15 => std_logic_vector(to_unsigned( 204, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 481 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 240, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 20, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 234, 8)),
10 => std_logic_vector(to_unsigned( 251, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 218, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 482 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 170, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 98, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 202, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 217, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 208, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 197, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 483 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 21, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 4, 8)),
7 => std_logic_vector(to_unsigned( 135, 8)),
8 => std_logic_vector(to_unsigned( 27, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 182, 8)),
14 => std_logic_vector(to_unsigned( 74, 8)),
15 => std_logic_vector(to_unsigned( 35, 8)),
16 => std_logic_vector(to_unsigned( 146, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 484 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 178, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 198, 8)),
6 => std_logic_vector(to_unsigned( 245, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 5, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 158, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 485 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 26, 8)),
3 => std_logic_vector(to_unsigned( 210, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 2, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 193, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 173, 8)),
14 => std_logic_vector(to_unsigned( 135, 8)),
15 => std_logic_vector(to_unsigned( 232, 8)),
16 => std_logic_vector(to_unsigned( 60, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 486 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 33, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 10, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 232, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 34, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 64, 8)),
14 => std_logic_vector(to_unsigned( 44, 8)),
15 => std_logic_vector(to_unsigned( 35, 8)),
16 => std_logic_vector(to_unsigned( 83, 8)),
17 => std_logic_vector(to_unsigned( 39, 8)),
18 => std_logic_vector(to_unsigned( 53, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 487 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 79, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 30, 8)),
5 => std_logic_vector(to_unsigned( 86, 8)),
6 => std_logic_vector(to_unsigned( 87, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 48, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 126, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011101
elsif count = 488 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 189, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 193, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 190, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 165, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 143, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 489 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 144, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 41, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 201, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 195, 8)),
11 => std_logic_vector(to_unsigned( 159, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 490 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 196, 8)),
3 => std_logic_vector(to_unsigned( 48, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 238, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 244, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 491 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 62, 8)),
3 => std_logic_vector(to_unsigned( 255, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 51, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 78, 8)),
12 => std_logic_vector(to_unsigned( 228, 8)),
13 => std_logic_vector(to_unsigned( 100, 8)),
14 => std_logic_vector(to_unsigned( 228, 8)),
15 => std_logic_vector(to_unsigned( 154, 8)),
16 => std_logic_vector(to_unsigned( 156, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 492 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 22, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 193, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 77, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 217, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 211, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 493 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 34, 8)),
2 => std_logic_vector(to_unsigned( 2, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 103, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 226, 8)),
9 => std_logic_vector(to_unsigned( 85, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 229, 8)),
14 => std_logic_vector(to_unsigned( 12, 8)),
15 => std_logic_vector(to_unsigned( 9, 8)),
16 => std_logic_vector(to_unsigned( 25, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 63, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110110
elsif count = 494 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 167, 8)),
2 => std_logic_vector(to_unsigned( 152, 8)),
3 => std_logic_vector(to_unsigned( 201, 8)),
4 => std_logic_vector(to_unsigned( 32, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 147, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 114, 8)),
10 => std_logic_vector(to_unsigned( 203, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 168, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 46, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 203, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 495 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 227, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 120, 8)),
9 => std_logic_vector(to_unsigned( 156, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 93, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 82, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 68, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 496 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 209, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 46, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 118, 8)),
10 => std_logic_vector(to_unsigned( 60, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 208, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 234, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 97, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 497 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 254, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 39, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 123, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 39, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 30, 8)),
13 => std_logic_vector(to_unsigned( 92, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 254, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 71, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 498 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 44, 8)),
3 => std_logic_vector(to_unsigned( 108, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 78, 8)),
6 => std_logic_vector(to_unsigned( 88, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 207, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 499 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 5, 8)),
4 => std_logic_vector(to_unsigned( 33, 8)),
5 => std_logic_vector(to_unsigned( 197, 8)),
6 => std_logic_vector(to_unsigned( 118, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 93, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 156, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 95, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 3, 8)),
15 => std_logic_vector(to_unsigned( 212, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 500 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 30, 8)),
3 => std_logic_vector(to_unsigned( 207, 8)),
4 => std_logic_vector(to_unsigned( 205, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 197, 8)),
7 => std_logic_vector(to_unsigned( 147, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 221, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 206, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 234, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 212, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 206, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 501 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 197, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 239, 8)),
5 => std_logic_vector(to_unsigned( 17, 8)),
6 => std_logic_vector(to_unsigned( 90, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 204, 8)),
9 => std_logic_vector(to_unsigned( 137, 8)),
10 => std_logic_vector(to_unsigned( 237, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 192, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 247, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 207, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 502 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 219, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 224, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 83, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 503 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 120, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 2, 8)),
8 => std_logic_vector(to_unsigned( 109, 8)),
9 => std_logic_vector(to_unsigned( 63, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 208, 8)),
14 => std_logic_vector(to_unsigned( 227, 8)),
15 => std_logic_vector(to_unsigned( 39, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 504 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 62, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 6, 8)),
8 => std_logic_vector(to_unsigned( 169, 8)),
9 => std_logic_vector(to_unsigned( 209, 8)),
10 => std_logic_vector(to_unsigned( 188, 8)),
11 => std_logic_vector(to_unsigned( 28, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 55, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 57, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 505 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 37, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 235, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 171, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 178, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 62, 8)),
13 => std_logic_vector(to_unsigned( 31, 8)),
14 => std_logic_vector(to_unsigned( 213, 8)),
15 => std_logic_vector(to_unsigned( 68, 8)),
16 => std_logic_vector(to_unsigned( 244, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 212, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 506 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 75, 8)),
2 => std_logic_vector(to_unsigned( 206, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 183, 8)),
5 => std_logic_vector(to_unsigned( 229, 8)),
6 => std_logic_vector(to_unsigned( 2, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 217, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 56, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 192, 8)),
13 => std_logic_vector(to_unsigned( 17, 8)),
14 => std_logic_vector(to_unsigned( 208, 8)),
15 => std_logic_vector(to_unsigned( 31, 8)),
16 => std_logic_vector(to_unsigned( 222, 8)),
17 => std_logic_vector(to_unsigned( 45, 8)),
18 => std_logic_vector(to_unsigned( 198, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 507 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 95, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 115, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 212, 8)),
8 => std_logic_vector(to_unsigned( 184, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 122, 8)),
11 => std_logic_vector(to_unsigned( 246, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 190, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 508 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 22, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 186, 8)),
12 => std_logic_vector(to_unsigned( 119, 8)),
13 => std_logic_vector(to_unsigned( 123, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 212, 8)),
16 => std_logic_vector(to_unsigned( 0, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 509 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 78, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 248, 8)),
6 => std_logic_vector(to_unsigned( 227, 8)),
7 => std_logic_vector(to_unsigned( 174, 8)),
8 => std_logic_vector(to_unsigned( 164, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 22, 8)),
13 => std_logic_vector(to_unsigned( 41, 8)),
14 => std_logic_vector(to_unsigned( 32, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 103, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 510 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 32, 8)),
2 => std_logic_vector(to_unsigned( 246, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 45, 8)),
7 => std_logic_vector(to_unsigned( 143, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 191, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 190, 8)),
12 => std_logic_vector(to_unsigned( 202, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 82, 8)),
15 => std_logic_vector(to_unsigned( 243, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 511 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 87, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 246, 8)),
9 => std_logic_vector(to_unsigned( 238, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 92, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 512 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 85, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 227, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 116, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 513 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 54, 8)),
2 => std_logic_vector(to_unsigned( 218, 8)),
3 => std_logic_vector(to_unsigned( 70, 8)),
4 => std_logic_vector(to_unsigned( 234, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 183, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 18, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 249, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 199, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011011
elsif count = 514 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 160, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 34, 8)),
10 => std_logic_vector(to_unsigned( 250, 8)),
11 => std_logic_vector(to_unsigned( 227, 8)),
12 => std_logic_vector(to_unsigned( 41, 8)),
13 => std_logic_vector(to_unsigned( 192, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 18, 8)),
16 => std_logic_vector(to_unsigned( 196, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 172, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00001111
elsif count = 515 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 147, 8)),
2 => std_logic_vector(to_unsigned( 141, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 85, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 120, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 58, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 119, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 516 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 166, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 50, 8)),
5 => std_logic_vector(to_unsigned( 63, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 42, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 34, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 230, 8)),
12 => std_logic_vector(to_unsigned( 38, 8)),
13 => std_logic_vector(to_unsigned( 29, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 170, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 517 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 224, 8)),
2 => std_logic_vector(to_unsigned( 76, 8)),
3 => std_logic_vector(to_unsigned( 129, 8)),
4 => std_logic_vector(to_unsigned( 187, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 108, 8)),
8 => std_logic_vector(to_unsigned( 228, 8)),
9 => std_logic_vector(to_unsigned( 90, 8)),
10 => std_logic_vector(to_unsigned( 210, 8)),
11 => std_logic_vector(to_unsigned( 246, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 32, 8)),
14 => std_logic_vector(to_unsigned( 240, 8)),
15 => std_logic_vector(to_unsigned( 103, 8)),
16 => std_logic_vector(to_unsigned( 223, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 198, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 518 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 210, 8)),
2 => std_logic_vector(to_unsigned( 188, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 247, 8)),
7 => std_logic_vector(to_unsigned( 217, 8)),
8 => std_logic_vector(to_unsigned( 36, 8)),
9 => std_logic_vector(to_unsigned( 45, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 193, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 208, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 187, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 203, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 519 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 8, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 59, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 29, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 25, 8)),
9 => std_logic_vector(to_unsigned( 86, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 213, 8)),
12 => std_logic_vector(to_unsigned( 32, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 7, 8)),
15 => std_logic_vector(to_unsigned( 238, 8)),
16 => std_logic_vector(to_unsigned( 50, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011011
elsif count = 520 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 184, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 9, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 83, 8)),
16 => std_logic_vector(to_unsigned( 214, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 57, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 521 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 54, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 7, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 47, 8)),
9 => std_logic_vector(to_unsigned( 84, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 186, 8)),
13 => std_logic_vector(to_unsigned( 50, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 18, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 522 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 216, 8)),
5 => std_logic_vector(to_unsigned( 159, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 94, 8)),
8 => std_logic_vector(to_unsigned( 93, 8)),
9 => std_logic_vector(to_unsigned( 14, 8)),
10 => std_logic_vector(to_unsigned( 137, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 31, 8)),
16 => std_logic_vector(to_unsigned( 7, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 523 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 64, 8)),
4 => std_logic_vector(to_unsigned( 214, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 198, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 206, 8)),
15 => std_logic_vector(to_unsigned( 78, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 524 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 82, 8)),
3 => std_logic_vector(to_unsigned( 20, 8)),
4 => std_logic_vector(to_unsigned( 102, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 202, 8)),
14 => std_logic_vector(to_unsigned( 73, 8)),
15 => std_logic_vector(to_unsigned( 55, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 525 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 224, 8)),
2 => std_logic_vector(to_unsigned( 83, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 213, 8)),
6 => std_logic_vector(to_unsigned( 72, 8)),
7 => std_logic_vector(to_unsigned( 235, 8)),
8 => std_logic_vector(to_unsigned( 94, 8)),
9 => std_logic_vector(to_unsigned( 182, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 131, 8)),
16 => std_logic_vector(to_unsigned( 50, 8)),
17 => std_logic_vector(to_unsigned( 205, 8)),
18 => std_logic_vector(to_unsigned( 106, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 526 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 91, 8)),
2 => std_logic_vector(to_unsigned( 64, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 250, 8)),
7 => std_logic_vector(to_unsigned( 250, 8)),
8 => std_logic_vector(to_unsigned( 40, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 23, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 63, 8)),
13 => std_logic_vector(to_unsigned( 45, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 8, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 61, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100011
elsif count = 527 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 1, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 173, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 63, 8)),
11 => std_logic_vector(to_unsigned( 186, 8)),
12 => std_logic_vector(to_unsigned( 162, 8)),
13 => std_logic_vector(to_unsigned( 183, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 528 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 231, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 189, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 130, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 51, 8)),
11 => std_logic_vector(to_unsigned( 218, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 529 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 237, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 154, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 53, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 107, 8)),
9 => std_logic_vector(to_unsigned( 22, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 21, 8)),
13 => std_logic_vector(to_unsigned( 56, 8)),
14 => std_logic_vector(to_unsigned( 32, 8)),
15 => std_logic_vector(to_unsigned( 254, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 530 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 96, 8)),
4 => std_logic_vector(to_unsigned( 36, 8)),
5 => std_logic_vector(to_unsigned( 40, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 73, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 531 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 129, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 230, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 94, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 26, 8)),
9 => std_logic_vector(to_unsigned( 177, 8)),
10 => std_logic_vector(to_unsigned( 15, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 39, 8)),
13 => std_logic_vector(to_unsigned( 212, 8)),
14 => std_logic_vector(to_unsigned( 52, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 63, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 51, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 532 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 255, 8)),
6 => std_logic_vector(to_unsigned( 210, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 37, 8)),
12 => std_logic_vector(to_unsigned( 70, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 533 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 68, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 233, 8)),
6 => std_logic_vector(to_unsigned( 15, 8)),
7 => std_logic_vector(to_unsigned( 252, 8)),
8 => std_logic_vector(to_unsigned( 218, 8)),
9 => std_logic_vector(to_unsigned( 126, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 136, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 47, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 215, 8)),
16 => std_logic_vector(to_unsigned( 28, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 158, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 534 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 229, 8)),
2 => std_logic_vector(to_unsigned( 121, 8)),
3 => std_logic_vector(to_unsigned( 231, 8)),
4 => std_logic_vector(to_unsigned( 119, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 254, 8)),
9 => std_logic_vector(to_unsigned( 231, 8)),
10 => std_logic_vector(to_unsigned( 119, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 23, 8)),
13 => std_logic_vector(to_unsigned( 225, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 535 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 130, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 205, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 195, 8)),
14 => std_logic_vector(to_unsigned( 1, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 105, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 536 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 242, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 192, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 208, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 189, 8)),
8 => std_logic_vector(to_unsigned( 37, 8)),
9 => std_logic_vector(to_unsigned( 144, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 139, 8)),
12 => std_logic_vector(to_unsigned( 79, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 243, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 537 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 241, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 202, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 234, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 197, 8)),
14 => std_logic_vector(to_unsigned( 218, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 164, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 538 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 8, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 60, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 71, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 126, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 539 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 139, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 112, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 14, 8)),
9 => std_logic_vector(to_unsigned( 78, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 13, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 69, 8)),
14 => std_logic_vector(to_unsigned( 69, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 53, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 43, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 540 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 13, 8)),
4 => std_logic_vector(to_unsigned( 16, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 238, 8)),
8 => std_logic_vector(to_unsigned( 185, 8)),
9 => std_logic_vector(to_unsigned( 112, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 31, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 541 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 176, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 39, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 235, 8)),
10 => std_logic_vector(to_unsigned( 173, 8)),
11 => std_logic_vector(to_unsigned( 48, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 105, 8)),
14 => std_logic_vector(to_unsigned( 181, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 190, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 542 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 147, 8)),
2 => std_logic_vector(to_unsigned( 195, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 141, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 225, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 543 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 94, 8)),
11 => std_logic_vector(to_unsigned( 75, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 228, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 544 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 91, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 114, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 50, 8)),
8 => std_logic_vector(to_unsigned( 75, 8)),
9 => std_logic_vector(to_unsigned( 118, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 545 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 131, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 78, 8)),
6 => std_logic_vector(to_unsigned( 228, 8)),
7 => std_logic_vector(to_unsigned( 183, 8)),
8 => std_logic_vector(to_unsigned( 165, 8)),
9 => std_logic_vector(to_unsigned( 134, 8)),
10 => std_logic_vector(to_unsigned( 180, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 218, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 546 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 127, 8)),
4 => std_logic_vector(to_unsigned( 129, 8)),
5 => std_logic_vector(to_unsigned( 96, 8)),
6 => std_logic_vector(to_unsigned( 200, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 46, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 238, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 234, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 547 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 194, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 89, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 131, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 160, 8)),
9 => std_logic_vector(to_unsigned( 152, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 179, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 144, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 548 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 73, 8)),
4 => std_logic_vector(to_unsigned( 106, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 166, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 231, 8)),
9 => std_logic_vector(to_unsigned( 23, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 98, 8)),
13 => std_logic_vector(to_unsigned( 219, 8)),
14 => std_logic_vector(to_unsigned( 13, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 164, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 549 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 203, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 171, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 230, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 188, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 182, 8)),
11 => std_logic_vector(to_unsigned( 224, 8)),
12 => std_logic_vector(to_unsigned( 173, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 191, 8)),
15 => std_logic_vector(to_unsigned( 100, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 200, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 550 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 224, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 213, 8)),
6 => std_logic_vector(to_unsigned( 199, 8)),
7 => std_logic_vector(to_unsigned( 208, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 187, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 66, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 61, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 551 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 41, 8)),
2 => std_logic_vector(to_unsigned( 193, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 184, 8)),
5 => std_logic_vector(to_unsigned( 47, 8)),
6 => std_logic_vector(to_unsigned( 115, 8)),
7 => std_logic_vector(to_unsigned( 242, 8)),
8 => std_logic_vector(to_unsigned( 251, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 33, 8)),
14 => std_logic_vector(to_unsigned( 119, 8)),
15 => std_logic_vector(to_unsigned( 36, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 42, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 552 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 85, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 197, 8)),
4 => std_logic_vector(to_unsigned( 66, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 22, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 228, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 36, 8)),
15 => std_logic_vector(to_unsigned( 194, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 553 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 249, 8)),
2 => std_logic_vector(to_unsigned( 82, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 235, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 15, 8)),
9 => std_logic_vector(to_unsigned( 51, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 219, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 195, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 554 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 232, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 220, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 96, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 74, 8)),
12 => std_logic_vector(to_unsigned( 223, 8)),
13 => std_logic_vector(to_unsigned( 66, 8)),
14 => std_logic_vector(to_unsigned( 215, 8)),
15 => std_logic_vector(to_unsigned( 52, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 555 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 177, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 207, 8)),
4 => std_logic_vector(to_unsigned( 13, 8)),
5 => std_logic_vector(to_unsigned( 158, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 231, 8)),
8 => std_logic_vector(to_unsigned( 44, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 139, 8)),
11 => std_logic_vector(to_unsigned( 112, 8)),
12 => std_logic_vector(to_unsigned( 239, 8)),
13 => std_logic_vector(to_unsigned( 222, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 91, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 556 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 37, 8)),
10 => std_logic_vector(to_unsigned( 159, 8)),
11 => std_logic_vector(to_unsigned( 156, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 33, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 557 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 128, 8)),
2 => std_logic_vector(to_unsigned( 177, 8)),
3 => std_logic_vector(to_unsigned( 149, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 141, 8)),
8 => std_logic_vector(to_unsigned( 7, 8)),
9 => std_logic_vector(to_unsigned( 176, 8)),
10 => std_logic_vector(to_unsigned( 189, 8)),
11 => std_logic_vector(to_unsigned( 213, 8)),
12 => std_logic_vector(to_unsigned( 12, 8)),
13 => std_logic_vector(to_unsigned( 138, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 9, 8)),
16 => std_logic_vector(to_unsigned( 225, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010011
elsif count = 558 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 1, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 169, 8)),
4 => std_logic_vector(to_unsigned( 204, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 197, 8)),
7 => std_logic_vector(to_unsigned( 229, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 220, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 80, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 559 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 150, 8)),
7 => std_logic_vector(to_unsigned( 209, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 184, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 0, 8)),
13 => std_logic_vector(to_unsigned( 155, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 560 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 227, 8)),
4 => std_logic_vector(to_unsigned( 217, 8)),
5 => std_logic_vector(to_unsigned( 224, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 191, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 157, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 182, 8)),
17 => std_logic_vector(to_unsigned( 155, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 561 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 29, 8)),
2 => std_logic_vector(to_unsigned( 188, 8)),
3 => std_logic_vector(to_unsigned( 106, 8)),
4 => std_logic_vector(to_unsigned( 49, 8)),
5 => std_logic_vector(to_unsigned( 134, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 75, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 35, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 153, 8)),
12 => std_logic_vector(to_unsigned( 96, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 562 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 39, 8)),
3 => std_logic_vector(to_unsigned( 13, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 51, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 177, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 74, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 237, 8)),
16 => std_logic_vector(to_unsigned( 119, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 563 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 247, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 109, 8)),
6 => std_logic_vector(to_unsigned( 217, 8)),
7 => std_logic_vector(to_unsigned( 83, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 227, 8)),
11 => std_logic_vector(to_unsigned( 221, 8)),
12 => std_logic_vector(to_unsigned( 151, 8)),
13 => std_logic_vector(to_unsigned( 133, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 71, 8)),
16 => std_logic_vector(to_unsigned( 175, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 564 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 71, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 173, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 137, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 128, 8)),
15 => std_logic_vector(to_unsigned( 16, 8)),
16 => std_logic_vector(to_unsigned( 252, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 565 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 29, 8)),
2 => std_logic_vector(to_unsigned( 41, 8)),
3 => std_logic_vector(to_unsigned( 62, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 21, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 252, 8)),
8 => std_logic_vector(to_unsigned( 234, 8)),
9 => std_logic_vector(to_unsigned( 39, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 14, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 44, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 49, 8)),
18 => std_logic_vector(to_unsigned( 197, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 566 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 152, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 18, 8)),
4 => std_logic_vector(to_unsigned( 59, 8)),
5 => std_logic_vector(to_unsigned( 41, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 17, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 84, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 9, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 6, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 68, 8)),
16 => std_logic_vector(to_unsigned( 118, 8)),
17 => std_logic_vector(to_unsigned( 45, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 567 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 45, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 207, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 217, 8)),
11 => std_logic_vector(to_unsigned( 153, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 209, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 223, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 209, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 568 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 52, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 112, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 112, 8)),
12 => std_logic_vector(to_unsigned( 201, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 20, 8)),
16 => std_logic_vector(to_unsigned( 26, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 569 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 96, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 214, 8)),
6 => std_logic_vector(to_unsigned( 209, 8)),
7 => std_logic_vector(to_unsigned( 85, 8)),
8 => std_logic_vector(to_unsigned( 211, 8)),
9 => std_logic_vector(to_unsigned( 60, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 177, 8)),
14 => std_logic_vector(to_unsigned( 147, 8)),
15 => std_logic_vector(to_unsigned( 6, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 570 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 154, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 166, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 94, 8)),
8 => std_logic_vector(to_unsigned( 130, 8)),
9 => std_logic_vector(to_unsigned( 190, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 134, 8)),
13 => std_logic_vector(to_unsigned( 205, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 571 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 11, 8)),
3 => std_logic_vector(to_unsigned( 110, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 116, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 112, 8)),
9 => std_logic_vector(to_unsigned( 10, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 66, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 67, 8)),
15 => std_logic_vector(to_unsigned( 238, 8)),
16 => std_logic_vector(to_unsigned( 238, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 91, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 572 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 128, 8)),
2 => std_logic_vector(to_unsigned( 141, 8)),
3 => std_logic_vector(to_unsigned( 224, 8)),
4 => std_logic_vector(to_unsigned( 40, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 112, 8)),
7 => std_logic_vector(to_unsigned( 19, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 137, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 87, 8)),
12 => std_logic_vector(to_unsigned( 29, 8)),
13 => std_logic_vector(to_unsigned( 65, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 231, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 573 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 18, 8)),
2 => std_logic_vector(to_unsigned( 16, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 18, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 38, 8)),
10 => std_logic_vector(to_unsigned( 184, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 126, 8)),
13 => std_logic_vector(to_unsigned( 39, 8)),
14 => std_logic_vector(to_unsigned( 177, 8)),
15 => std_logic_vector(to_unsigned( 253, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 181, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 574 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 191, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 141, 8)),
6 => std_logic_vector(to_unsigned( 229, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 240, 8)),
9 => std_logic_vector(to_unsigned( 80, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 210, 8)),
13 => std_logic_vector(to_unsigned( 15, 8)),
14 => std_logic_vector(to_unsigned( 67, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 203, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 177, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 575 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 229, 8)),
2 => std_logic_vector(to_unsigned( 201, 8)),
3 => std_logic_vector(to_unsigned( 219, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 185, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 89, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 141, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 576 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 218, 8)),
2 => std_logic_vector(to_unsigned( 64, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 224, 8)),
6 => std_logic_vector(to_unsigned( 70, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 52, 8)),
9 => std_logic_vector(to_unsigned( 54, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 226, 8)),
13 => std_logic_vector(to_unsigned( 26, 8)),
14 => std_logic_vector(to_unsigned( 51, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 577 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 99, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 78, 8)),
4 => std_logic_vector(to_unsigned( 10, 8)),
5 => std_logic_vector(to_unsigned( 32, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 86, 8)),
8 => std_logic_vector(to_unsigned( 16, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 94, 8)),
11 => std_logic_vector(to_unsigned( 54, 8)),
12 => std_logic_vector(to_unsigned( 34, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 243, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 75, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 578 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 91, 8)),
5 => std_logic_vector(to_unsigned( 165, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 2, 8)),
14 => std_logic_vector(to_unsigned( 178, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 579 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 143, 8)),
2 => std_logic_vector(to_unsigned( 151, 8)),
3 => std_logic_vector(to_unsigned( 48, 8)),
4 => std_logic_vector(to_unsigned( 2, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 20, 8)),
9 => std_logic_vector(to_unsigned( 93, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 33, 8)),
13 => std_logic_vector(to_unsigned( 13, 8)),
14 => std_logic_vector(to_unsigned( 255, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010101
elsif count = 580 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 10, 8)),
6 => std_logic_vector(to_unsigned( 241, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 77, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 83, 8)),
13 => std_logic_vector(to_unsigned( 155, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 61, 8)),
16 => std_logic_vector(to_unsigned( 252, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 581 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 2, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 30, 8)),
6 => std_logic_vector(to_unsigned( 236, 8)),
7 => std_logic_vector(to_unsigned( 102, 8)),
8 => std_logic_vector(to_unsigned( 42, 8)),
9 => std_logic_vector(to_unsigned( 80, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 119, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 582 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 96, 8)),
5 => std_logic_vector(to_unsigned( 8, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 2, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 161, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010011
elsif count = 583 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 167, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 225, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 58, 8)),
8 => std_logic_vector(to_unsigned( 120, 8)),
9 => std_logic_vector(to_unsigned( 63, 8)),
10 => std_logic_vector(to_unsigned( 115, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 71, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 57, 8)),
16 => std_logic_vector(to_unsigned( 121, 8)),
17 => std_logic_vector(to_unsigned( 50, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 584 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 158, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 201, 8)),
5 => std_logic_vector(to_unsigned( 159, 8)),
6 => std_logic_vector(to_unsigned( 213, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 217, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 92, 8)),
13 => std_logic_vector(to_unsigned( 154, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 5, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 186, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 585 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 166, 8)),
2 => std_logic_vector(to_unsigned( 217, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 233, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 226, 8)),
9 => std_logic_vector(to_unsigned( 230, 8)),
10 => std_logic_vector(to_unsigned( 185, 8)),
11 => std_logic_vector(to_unsigned( 144, 8)),
12 => std_logic_vector(to_unsigned( 255, 8)),
13 => std_logic_vector(to_unsigned( 170, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 197, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 586 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 132, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 204, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 19, 8)),
7 => std_logic_vector(to_unsigned( 44, 8)),
8 => std_logic_vector(to_unsigned( 140, 8)),
9 => std_logic_vector(to_unsigned( 53, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 95, 8)),
13 => std_logic_vector(to_unsigned( 200, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010011
elsif count = 587 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 241, 8)),
5 => std_logic_vector(to_unsigned( 171, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 204, 8)),
8 => std_logic_vector(to_unsigned( 17, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 0, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 3, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 53, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 588 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 183, 8)),
3 => std_logic_vector(to_unsigned( 123, 8)),
4 => std_logic_vector(to_unsigned( 223, 8)),
5 => std_logic_vector(to_unsigned( 109, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 220, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 174, 8)),
11 => std_logic_vector(to_unsigned( 244, 8)),
12 => std_logic_vector(to_unsigned( 19, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 9, 8)),
15 => std_logic_vector(to_unsigned( 127, 8)),
16 => std_logic_vector(to_unsigned( 219, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 198, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 589 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 47, 8)),
5 => std_logic_vector(to_unsigned( 76, 8)),
6 => std_logic_vector(to_unsigned( 37, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 246, 8)),
10 => std_logic_vector(to_unsigned( 214, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 39, 8)),
13 => std_logic_vector(to_unsigned( 59, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 234, 8)),
16 => std_logic_vector(to_unsigned( 237, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 590 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 24, 8)),
2 => std_logic_vector(to_unsigned( 3, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 35, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 243, 8)),
15 => std_logic_vector(to_unsigned( 38, 8)),
16 => std_logic_vector(to_unsigned( 20, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 591 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 228, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 222, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 95, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 250, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 201, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 18, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100100
elsif count = 592 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 58, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 86, 8)),
6 => std_logic_vector(to_unsigned( 168, 8)),
7 => std_logic_vector(to_unsigned( 50, 8)),
8 => std_logic_vector(to_unsigned( 35, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 130, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 51, 8)),
13 => std_logic_vector(to_unsigned( 179, 8)),
14 => std_logic_vector(to_unsigned( 131, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 75, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 593 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 81, 8)),
3 => std_logic_vector(to_unsigned( 234, 8)),
4 => std_logic_vector(to_unsigned( 226, 8)),
5 => std_logic_vector(to_unsigned( 254, 8)),
6 => std_logic_vector(to_unsigned( 235, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 39, 8)),
10 => std_logic_vector(to_unsigned( 125, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 202, 8)),
15 => std_logic_vector(to_unsigned( 187, 8)),
16 => std_logic_vector(to_unsigned( 198, 8)),
17 => std_logic_vector(to_unsigned( 219, 8)),
18 => std_logic_vector(to_unsigned( 211, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 594 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 61, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 227, 8)),
6 => std_logic_vector(to_unsigned( 95, 8)),
7 => std_logic_vector(to_unsigned( 181, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 191, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 152, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 184, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 595 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 38, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 181, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 217, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 596 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 67, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 12, 8)),
6 => std_logic_vector(to_unsigned( 169, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 51, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 105, 8)),
15 => std_logic_vector(to_unsigned( 24, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 597 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 83, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 171, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 93, 8)),
6 => std_logic_vector(to_unsigned( 26, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 93, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 31, 8)),
14 => std_logic_vector(to_unsigned( 131, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 170, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 598 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 211, 8)),
2 => std_logic_vector(to_unsigned( 11, 8)),
3 => std_logic_vector(to_unsigned( 217, 8)),
4 => std_logic_vector(to_unsigned( 45, 8)),
5 => std_logic_vector(to_unsigned( 231, 8)),
6 => std_logic_vector(to_unsigned( 31, 8)),
7 => std_logic_vector(to_unsigned( 150, 8)),
8 => std_logic_vector(to_unsigned( 81, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 7, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 29, 8)),
13 => std_logic_vector(to_unsigned( 200, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 254, 8)),
17 => std_logic_vector(to_unsigned( 200, 8)),
18 => std_logic_vector(to_unsigned( 31, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 599 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 18, 8)),
2 => std_logic_vector(to_unsigned( 48, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 234, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 58, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001110
elsif count = 600 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 68, 8)),
3 => std_logic_vector(to_unsigned( 112, 8)),
4 => std_logic_vector(to_unsigned( 53, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 209, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 193, 8)),
9 => std_logic_vector(to_unsigned( 99, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 128, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 601 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 68, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 144, 8)),
9 => std_logic_vector(to_unsigned( 218, 8)),
10 => std_logic_vector(to_unsigned( 59, 8)),
11 => std_logic_vector(to_unsigned( 43, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 230, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 249, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 602 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 39, 8)),
7 => std_logic_vector(to_unsigned( 50, 8)),
8 => std_logic_vector(to_unsigned( 221, 8)),
9 => std_logic_vector(to_unsigned( 100, 8)),
10 => std_logic_vector(to_unsigned( 46, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 78, 8)),
16 => std_logic_vector(to_unsigned( 68, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 603 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 193, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 231, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 200, 8)),
11 => std_logic_vector(to_unsigned( 252, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 102, 8)),
14 => std_logic_vector(to_unsigned( 211, 8)),
15 => std_logic_vector(to_unsigned( 230, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 75, 8)),
18 => std_logic_vector(to_unsigned( 214, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 604 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 83, 8)),
7 => std_logic_vector(to_unsigned( 161, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 136, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 203, 8)),
12 => std_logic_vector(to_unsigned( 47, 8)),
13 => std_logic_vector(to_unsigned( 201, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 191, 8)),
16 => std_logic_vector(to_unsigned( 9, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 605 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 22, 8)),
2 => std_logic_vector(to_unsigned( 38, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 202, 8)),
6 => std_logic_vector(to_unsigned( 58, 8)),
7 => std_logic_vector(to_unsigned( 174, 8)),
8 => std_logic_vector(to_unsigned( 30, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 211, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 606 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 40, 8)),
2 => std_logic_vector(to_unsigned( 187, 8)),
3 => std_logic_vector(to_unsigned( 81, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 24, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 188, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 246, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 168, 8)),
16 => std_logic_vector(to_unsigned( 153, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110010
elsif count = 607 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 182, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 154, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 182, 8)),
7 => std_logic_vector(to_unsigned( 208, 8)),
8 => std_logic_vector(to_unsigned( 131, 8)),
9 => std_logic_vector(to_unsigned( 199, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 177, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 608 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 164, 8)),
5 => std_logic_vector(to_unsigned( 183, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 176, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 181, 8)),
10 => std_logic_vector(to_unsigned( 96, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 205, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 609 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 125, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 88, 8)),
6 => std_logic_vector(to_unsigned( 115, 8)),
7 => std_logic_vector(to_unsigned( 34, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 80, 8)),
12 => std_logic_vector(to_unsigned( 193, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 195, 8)),
15 => std_logic_vector(to_unsigned( 237, 8)),
16 => std_logic_vector(to_unsigned( 205, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 610 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 249, 8)),
3 => std_logic_vector(to_unsigned( 235, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 103, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 208, 8)),
8 => std_logic_vector(to_unsigned( 46, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 145, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 119, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 130, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 611 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 71, 8)),
3 => std_logic_vector(to_unsigned( 231, 8)),
4 => std_logic_vector(to_unsigned( 73, 8)),
5 => std_logic_vector(to_unsigned( 93, 8)),
6 => std_logic_vector(to_unsigned( 98, 8)),
7 => std_logic_vector(to_unsigned( 206, 8)),
8 => std_logic_vector(to_unsigned( 112, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 169, 8)),
14 => std_logic_vector(to_unsigned( 71, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 47, 8)),
17 => std_logic_vector(to_unsigned( 199, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 612 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 237, 8)),
5 => std_logic_vector(to_unsigned( 52, 8)),
6 => std_logic_vector(to_unsigned( 4, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 139, 8)),
11 => std_logic_vector(to_unsigned( 51, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 140, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011000
elsif count = 613 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 221, 8)),
2 => std_logic_vector(to_unsigned( 10, 8)),
3 => std_logic_vector(to_unsigned( 185, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 198, 8)),
8 => std_logic_vector(to_unsigned( 151, 8)),
9 => std_logic_vector(to_unsigned( 206, 8)),
10 => std_logic_vector(to_unsigned( 215, 8)),
11 => std_logic_vector(to_unsigned( 232, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 154, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 187, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 614 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 162, 8)),
2 => std_logic_vector(to_unsigned( 60, 8)),
3 => std_logic_vector(to_unsigned( 233, 8)),
4 => std_logic_vector(to_unsigned( 22, 8)),
5 => std_logic_vector(to_unsigned( 183, 8)),
6 => std_logic_vector(to_unsigned( 17, 8)),
7 => std_logic_vector(to_unsigned( 222, 8)),
8 => std_logic_vector(to_unsigned( 143, 8)),
9 => std_logic_vector(to_unsigned( 160, 8)),
10 => std_logic_vector(to_unsigned( 30, 8)),
11 => std_logic_vector(to_unsigned( 243, 8)),
12 => std_logic_vector(to_unsigned( 43, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 204, 8)),
16 => std_logic_vector(to_unsigned( 197, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 44, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 615 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 95, 8)),
2 => std_logic_vector(to_unsigned( 155, 8)),
3 => std_logic_vector(to_unsigned( 51, 8)),
4 => std_logic_vector(to_unsigned( 99, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 13, 8)),
7 => std_logic_vector(to_unsigned( 245, 8)),
8 => std_logic_vector(to_unsigned( 196, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 107, 8)),
11 => std_logic_vector(to_unsigned( 120, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 227, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 123, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 616 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 24, 8)),
5 => std_logic_vector(to_unsigned( 147, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 63, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 207, 8)),
12 => std_logic_vector(to_unsigned( 116, 8)),
13 => std_logic_vector(to_unsigned( 158, 8)),
14 => std_logic_vector(to_unsigned( 163, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 195, 8)),
17 => std_logic_vector(to_unsigned( 206, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 617 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 125, 8)),
3 => std_logic_vector(to_unsigned( 35, 8)),
4 => std_logic_vector(to_unsigned( 79, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 105, 8)),
7 => std_logic_vector(to_unsigned( 152, 8)),
8 => std_logic_vector(to_unsigned( 6, 8)),
9 => std_logic_vector(to_unsigned( 244, 8)),
10 => std_logic_vector(to_unsigned( 206, 8)),
11 => std_logic_vector(to_unsigned( 49, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 254, 8)),
14 => std_logic_vector(to_unsigned( 165, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 52, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 618 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 136, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 216, 8)),
5 => std_logic_vector(to_unsigned( 53, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 229, 8)),
11 => std_logic_vector(to_unsigned( 5, 8)),
12 => std_logic_vector(to_unsigned( 5, 8)),
13 => std_logic_vector(to_unsigned( 2, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 21, 8)),
16 => std_logic_vector(to_unsigned( 138, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 619 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 169, 8)),
3 => std_logic_vector(to_unsigned( 92, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 63, 8)),
6 => std_logic_vector(to_unsigned( 173, 8)),
7 => std_logic_vector(to_unsigned( 3, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 0, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 248, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 167, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 118, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 620 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 203, 8)),
2 => std_logic_vector(to_unsigned( 45, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 7, 8)),
5 => std_logic_vector(to_unsigned( 253, 8)),
6 => std_logic_vector(to_unsigned( 114, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 155, 8)),
10 => std_logic_vector(to_unsigned( 166, 8)),
11 => std_logic_vector(to_unsigned( 196, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 193, 8)),
16 => std_logic_vector(to_unsigned( 30, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 621 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 250, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 226, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 228, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 64, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 142, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 143, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 622 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 213, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 26, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 52, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 130, 8)),
15 => std_logic_vector(to_unsigned( 12, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 153, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110101
elsif count = 623 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 16, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 18, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 120, 8)),
12 => std_logic_vector(to_unsigned( 73, 8)),
13 => std_logic_vector(to_unsigned( 25, 8)),
14 => std_logic_vector(to_unsigned( 83, 8)),
15 => std_logic_vector(to_unsigned( 35, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 624 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 150, 8)),
2 => std_logic_vector(to_unsigned( 153, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 103, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 196, 8)),
8 => std_logic_vector(to_unsigned( 60, 8)),
9 => std_logic_vector(to_unsigned( 23, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 157, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 195, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 625 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 31, 8)),
8 => std_logic_vector(to_unsigned( 189, 8)),
9 => std_logic_vector(to_unsigned( 177, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 198, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 145, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 626 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 243, 8)),
3 => std_logic_vector(to_unsigned( 113, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 173, 8)),
6 => std_logic_vector(to_unsigned( 25, 8)),
7 => std_logic_vector(to_unsigned( 19, 8)),
8 => std_logic_vector(to_unsigned( 0, 8)),
9 => std_logic_vector(to_unsigned( 163, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 159, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 236, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 59, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110100
elsif count = 627 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 61, 8)),
2 => std_logic_vector(to_unsigned( 29, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 193, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 30, 8)),
7 => std_logic_vector(to_unsigned( 203, 8)),
8 => std_logic_vector(to_unsigned( 166, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 20, 8)),
11 => std_logic_vector(to_unsigned( 190, 8)),
12 => std_logic_vector(to_unsigned( 233, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 214, 8)),
15 => std_logic_vector(to_unsigned( 240, 8)),
16 => std_logic_vector(to_unsigned( 203, 8)),
17 => std_logic_vector(to_unsigned( 203, 8)),
18 => std_logic_vector(to_unsigned( 206, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101010
elsif count = 628 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 49, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 30, 8)),
6 => std_logic_vector(to_unsigned( 159, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 247, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 85, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 135, 8)),
14 => std_logic_vector(to_unsigned( 182, 8)),
15 => std_logic_vector(to_unsigned( 128, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 629 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 59, 8)),
4 => std_logic_vector(to_unsigned( 245, 8)),
5 => std_logic_vector(to_unsigned( 133, 8)),
6 => std_logic_vector(to_unsigned( 38, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 188, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 51, 8)),
13 => std_logic_vector(to_unsigned( 202, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 227, 8)),
16 => std_logic_vector(to_unsigned( 242, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 630 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 71, 8)),
2 => std_logic_vector(to_unsigned( 122, 8)),
3 => std_logic_vector(to_unsigned( 61, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 152, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 82, 8)),
11 => std_logic_vector(to_unsigned( 198, 8)),
12 => std_logic_vector(to_unsigned( 131, 8)),
13 => std_logic_vector(to_unsigned( 97, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 72, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 631 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 103, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 16, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 56, 8)),
10 => std_logic_vector(to_unsigned( 155, 8)),
11 => std_logic_vector(to_unsigned( 13, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 81, 8)),
16 => std_logic_vector(to_unsigned( 80, 8)),
17 => std_logic_vector(to_unsigned( 58, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 632 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 72, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 66, 8)),
5 => std_logic_vector(to_unsigned( 76, 8)),
6 => std_logic_vector(to_unsigned( 50, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 31, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 191, 8)),
13 => std_logic_vector(to_unsigned( 64, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 251, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 633 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 144, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 234, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 69, 8)),
15 => std_logic_vector(to_unsigned( 90, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 634 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 92, 8)),
3 => std_logic_vector(to_unsigned( 245, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 146, 8)),
6 => std_logic_vector(to_unsigned( 16, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 221, 8)),
10 => std_logic_vector(to_unsigned( 124, 8)),
11 => std_logic_vector(to_unsigned( 63, 8)),
12 => std_logic_vector(to_unsigned( 51, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 635 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 211, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 79, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 77, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 64, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 74, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001110
elsif count = 636 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 147, 8)),
2 => std_logic_vector(to_unsigned( 136, 8)),
3 => std_logic_vector(to_unsigned( 238, 8)),
4 => std_logic_vector(to_unsigned( 63, 8)),
5 => std_logic_vector(to_unsigned( 68, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 213, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 209, 8)),
13 => std_logic_vector(to_unsigned( 28, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 196, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 637 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 246, 8)),
3 => std_logic_vector(to_unsigned( 9, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 225, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 165, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 243, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 64, 8)),
18 => std_logic_vector(to_unsigned( 132, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 638 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 132, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 148, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 136, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 5, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 639 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 124, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 182, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 120, 8)),
15 => std_logic_vector(to_unsigned( 22, 8)),
16 => std_logic_vector(to_unsigned( 181, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 161, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 640 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 249, 8)),
2 => std_logic_vector(to_unsigned( 151, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 97, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 199, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 62, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 15, 8)),
12 => std_logic_vector(to_unsigned( 173, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 111, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001010
elsif count = 641 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 186, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 166, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 15, 8)),
7 => std_logic_vector(to_unsigned( 189, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 97, 8)),
15 => std_logic_vector(to_unsigned( 205, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 642 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 80, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 233, 8)),
4 => std_logic_vector(to_unsigned( 187, 8)),
5 => std_logic_vector(to_unsigned( 28, 8)),
6 => std_logic_vector(to_unsigned( 70, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 109, 8)),
10 => std_logic_vector(to_unsigned( 166, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 72, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 643 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 223, 8)),
3 => std_logic_vector(to_unsigned( 103, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 174, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 193, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 644 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 136, 8)),
3 => std_logic_vector(to_unsigned( 172, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 144, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 250, 8)),
13 => std_logic_vector(to_unsigned( 2, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 645 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 88, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 72, 8)),
5 => std_logic_vector(to_unsigned( 116, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 111, 8)),
10 => std_logic_vector(to_unsigned( 253, 8)),
11 => std_logic_vector(to_unsigned( 45, 8)),
12 => std_logic_vector(to_unsigned( 38, 8)),
13 => std_logic_vector(to_unsigned( 21, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 646 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 62, 8)),
4 => std_logic_vector(to_unsigned( 166, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 45, 8)),
8 => std_logic_vector(to_unsigned( 250, 8)),
9 => std_logic_vector(to_unsigned( 179, 8)),
10 => std_logic_vector(to_unsigned( 8, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 33, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 187, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 166, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 647 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 129, 8)),
2 => std_logic_vector(to_unsigned( 212, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 76, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 83, 8)),
7 => std_logic_vector(to_unsigned( 154, 8)),
8 => std_logic_vector(to_unsigned( 36, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 36, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 69, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 61, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 648 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 91, 8)),
4 => std_logic_vector(to_unsigned( 238, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 195, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 21, 8)),
11 => std_logic_vector(to_unsigned( 44, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 165, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 649 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 70, 8)),
4 => std_logic_vector(to_unsigned( 168, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 41, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 29, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 650 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 225, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 80, 8)),
7 => std_logic_vector(to_unsigned( 222, 8)),
8 => std_logic_vector(to_unsigned( 38, 8)),
9 => std_logic_vector(to_unsigned( 202, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 231, 8)),
14 => std_logic_vector(to_unsigned( 54, 8)),
15 => std_logic_vector(to_unsigned( 235, 8)),
16 => std_logic_vector(to_unsigned( 58, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 651 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 185, 8)),
2 => std_logic_vector(to_unsigned( 63, 8)),
3 => std_logic_vector(to_unsigned( 14, 8)),
4 => std_logic_vector(to_unsigned( 211, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 193, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 181, 8)),
10 => std_logic_vector(to_unsigned( 179, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 249, 8)),
14 => std_logic_vector(to_unsigned( 113, 8)),
15 => std_logic_vector(to_unsigned( 251, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 205, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 652 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 198, 8)),
3 => std_logic_vector(to_unsigned( 229, 8)),
4 => std_logic_vector(to_unsigned( 16, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 37, 8)),
9 => std_logic_vector(to_unsigned( 254, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 198, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 77, 8)),
15 => std_logic_vector(to_unsigned( 181, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100100
elsif count = 653 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 157, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 5, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 221, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 225, 8)),
8 => std_logic_vector(to_unsigned( 85, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 87, 8)),
11 => std_logic_vector(to_unsigned( 246, 8)),
12 => std_logic_vector(to_unsigned( 3, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 208, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 654 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 7, 8)),
3 => std_logic_vector(to_unsigned( 67, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 20, 8)),
8 => std_logic_vector(to_unsigned( 78, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 122, 8)),
11 => std_logic_vector(to_unsigned( 101, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 132, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 75, 8)),
18 => std_logic_vector(to_unsigned( 81, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 655 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 124, 8)),
8 => std_logic_vector(to_unsigned( 81, 8)),
9 => std_logic_vector(to_unsigned( 138, 8)),
10 => std_logic_vector(to_unsigned( 95, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 184, 8)),
13 => std_logic_vector(to_unsigned( 46, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 153, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 656 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 118, 8)),
3 => std_logic_vector(to_unsigned( 243, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 146, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 115, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 167, 8)),
16 => std_logic_vector(to_unsigned( 33, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 657 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 250, 8)),
4 => std_logic_vector(to_unsigned( 238, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 230, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 79, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 18, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 658 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 160, 8)),
3 => std_logic_vector(to_unsigned( 14, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 34, 8)),
7 => std_logic_vector(to_unsigned( 148, 8)),
8 => std_logic_vector(to_unsigned( 225, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 58, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 86, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 78, 8)),
15 => std_logic_vector(to_unsigned( 54, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 659 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 78, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 173, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 206, 8)),
12 => std_logic_vector(to_unsigned( 6, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 79, 8)),
15 => std_logic_vector(to_unsigned( 99, 8)),
16 => std_logic_vector(to_unsigned( 155, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 660 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 74, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 243, 8)),
4 => std_logic_vector(to_unsigned( 118, 8)),
5 => std_logic_vector(to_unsigned( 203, 8)),
6 => std_logic_vector(to_unsigned( 173, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 37, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 176, 8)),
11 => std_logic_vector(to_unsigned( 153, 8)),
12 => std_logic_vector(to_unsigned( 135, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 61, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001001
elsif count = 661 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 45, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 93, 8)),
9 => std_logic_vector(to_unsigned( 134, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 5, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 187, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 41, 8)),
17 => std_logic_vector(to_unsigned( 150, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 662 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 6, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 125, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 250, 8)),
9 => std_logic_vector(to_unsigned( 72, 8)),
10 => std_logic_vector(to_unsigned( 124, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 42, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 226, 8)),
16 => std_logic_vector(to_unsigned( 52, 8)),
17 => std_logic_vector(to_unsigned( 102, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 663 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 242, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 39, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 56, 8)),
10 => std_logic_vector(to_unsigned( 71, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 192, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 53, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100101
elsif count = 664 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 34, 8)),
3 => std_logic_vector(to_unsigned( 197, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 73, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 126, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 215, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 52, 8)),
13 => std_logic_vector(to_unsigned( 137, 8)),
14 => std_logic_vector(to_unsigned( 56, 8)),
15 => std_logic_vector(to_unsigned( 230, 8)),
16 => std_logic_vector(to_unsigned( 132, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 86, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 665 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 134, 8)),
5 => std_logic_vector(to_unsigned( 146, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 96, 8)),
13 => std_logic_vector(to_unsigned( 202, 8)),
14 => std_logic_vector(to_unsigned( 105, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 666 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 2, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 242, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 221, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 192, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 229, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 114, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 667 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 129, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 61, 8)),
5 => std_logic_vector(to_unsigned( 101, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 67, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 152, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 168, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 668 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 166, 8)),
2 => std_logic_vector(to_unsigned( 88, 8)),
3 => std_logic_vector(to_unsigned( 37, 8)),
4 => std_logic_vector(to_unsigned( 7, 8)),
5 => std_logic_vector(to_unsigned( 204, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 176, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 213, 8)),
10 => std_logic_vector(to_unsigned( 135, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 169, 8)),
13 => std_logic_vector(to_unsigned( 184, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 200, 8)),
18 => std_logic_vector(to_unsigned( 154, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111100
elsif count = 669 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 51, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 223, 8)),
4 => std_logic_vector(to_unsigned( 125, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 237, 8)),
7 => std_logic_vector(to_unsigned( 84, 8)),
8 => std_logic_vector(to_unsigned( 161, 8)),
9 => std_logic_vector(to_unsigned( 250, 8)),
10 => std_logic_vector(to_unsigned( 215, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 115, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 670 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 236, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 163, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 34, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 138, 8)),
16 => std_logic_vector(to_unsigned( 18, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 60, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111100
elsif count = 671 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 60, 8)),
3 => std_logic_vector(to_unsigned( 17, 8)),
4 => std_logic_vector(to_unsigned( 13, 8)),
5 => std_logic_vector(to_unsigned( 23, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 239, 8)),
8 => std_logic_vector(to_unsigned( 240, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 36, 8)),
12 => std_logic_vector(to_unsigned( 132, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 136, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 672 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 229, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 236, 8)),
6 => std_logic_vector(to_unsigned( 21, 8)),
7 => std_logic_vector(to_unsigned( 89, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 227, 8)),
10 => std_logic_vector(to_unsigned( 39, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 253, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 226, 8)),
15 => std_logic_vector(to_unsigned( 46, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 673 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 146, 8)),
3 => std_logic_vector(to_unsigned( 151, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 206, 8)),
12 => std_logic_vector(to_unsigned( 23, 8)),
13 => std_logic_vector(to_unsigned( 42, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 33, 8)),
16 => std_logic_vector(to_unsigned( 49, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 49, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 674 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 152, 8)),
2 => std_logic_vector(to_unsigned( 131, 8)),
3 => std_logic_vector(to_unsigned( 124, 8)),
4 => std_logic_vector(to_unsigned( 159, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 67, 8)),
8 => std_logic_vector(to_unsigned( 86, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 44, 8)),
14 => std_logic_vector(to_unsigned( 245, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 675 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 118, 8)),
2 => std_logic_vector(to_unsigned( 187, 8)),
3 => std_logic_vector(to_unsigned( 59, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 212, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 81, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 29, 8)),
12 => std_logic_vector(to_unsigned( 23, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 195, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 676 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 80, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 169, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 36, 8)),
10 => std_logic_vector(to_unsigned( 214, 8)),
11 => std_logic_vector(to_unsigned( 96, 8)),
12 => std_logic_vector(to_unsigned( 166, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 125, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 677 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 230, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 206, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 9, 8)),
9 => std_logic_vector(to_unsigned( 190, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 35, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 227, 8)),
16 => std_logic_vector(to_unsigned( 209, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 200, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110110
elsif count = 678 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 79, 8)),
4 => std_logic_vector(to_unsigned( 79, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 164, 8)),
7 => std_logic_vector(to_unsigned( 231, 8)),
8 => std_logic_vector(to_unsigned( 230, 8)),
9 => std_logic_vector(to_unsigned( 19, 8)),
10 => std_logic_vector(to_unsigned( 218, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 679 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 3, 8)),
2 => std_logic_vector(to_unsigned( 64, 8)),
3 => std_logic_vector(to_unsigned( 23, 8)),
4 => std_logic_vector(to_unsigned( 102, 8)),
5 => std_logic_vector(to_unsigned( 40, 8)),
6 => std_logic_vector(to_unsigned( 27, 8)),
7 => std_logic_vector(to_unsigned( 101, 8)),
8 => std_logic_vector(to_unsigned( 56, 8)),
9 => std_logic_vector(to_unsigned( 56, 8)),
10 => std_logic_vector(to_unsigned( 11, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 4, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 210, 8)),
16 => std_logic_vector(to_unsigned( 19, 8)),
17 => std_logic_vector(to_unsigned( 56, 8)),
18 => std_logic_vector(to_unsigned( 67, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 680 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 91, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 91, 8)),
4 => std_logic_vector(to_unsigned( 51, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 254, 8)),
8 => std_logic_vector(to_unsigned( 223, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 56, 8)),
12 => std_logic_vector(to_unsigned( 100, 8)),
13 => std_logic_vector(to_unsigned( 195, 8)),
14 => std_logic_vector(to_unsigned( 83, 8)),
15 => std_logic_vector(to_unsigned( 96, 8)),
16 => std_logic_vector(to_unsigned( 255, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 681 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 54, 8)),
3 => std_logic_vector(to_unsigned( 3, 8)),
4 => std_logic_vector(to_unsigned( 254, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 50, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 10, 8)),
9 => std_logic_vector(to_unsigned( 203, 8)),
10 => std_logic_vector(to_unsigned( 59, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 221, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 251, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 53, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111100
elsif count = 682 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 200, 8)),
2 => std_logic_vector(to_unsigned( 45, 8)),
3 => std_logic_vector(to_unsigned( 229, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 228, 8)),
6 => std_logic_vector(to_unsigned( 53, 8)),
7 => std_logic_vector(to_unsigned( 73, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 229, 8)),
10 => std_logic_vector(to_unsigned( 14, 8)),
11 => std_logic_vector(to_unsigned( 63, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 223, 8)),
14 => std_logic_vector(to_unsigned( 8, 8)),
15 => std_logic_vector(to_unsigned( 220, 8)),
16 => std_logic_vector(to_unsigned( 5, 8)),
17 => std_logic_vector(to_unsigned( 218, 8)),
18 => std_logic_vector(to_unsigned( 33, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 683 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 104, 8)),
2 => std_logic_vector(to_unsigned( 201, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 255, 8)),
7 => std_logic_vector(to_unsigned( 222, 8)),
8 => std_logic_vector(to_unsigned( 230, 8)),
9 => std_logic_vector(to_unsigned( 205, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 214, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 154, 8)),
14 => std_logic_vector(to_unsigned( 47, 8)),
15 => std_logic_vector(to_unsigned( 154, 8)),
16 => std_logic_vector(to_unsigned( 98, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110010
elsif count = 684 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 49, 8)),
4 => std_logic_vector(to_unsigned( 219, 8)),
5 => std_logic_vector(to_unsigned( 91, 8)),
6 => std_logic_vector(to_unsigned( 204, 8)),
7 => std_logic_vector(to_unsigned( 46, 8)),
8 => std_logic_vector(to_unsigned( 118, 8)),
9 => std_logic_vector(to_unsigned( 130, 8)),
10 => std_logic_vector(to_unsigned( 128, 8)),
11 => std_logic_vector(to_unsigned( 44, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 93, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111001
elsif count = 685 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 70, 8)),
4 => std_logic_vector(to_unsigned( 215, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 98, 8)),
8 => std_logic_vector(to_unsigned( 140, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 20, 8)),
16 => std_logic_vector(to_unsigned( 222, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 686 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 25, 8)),
3 => std_logic_vector(to_unsigned( 43, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 17, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 24, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 213, 8)),
12 => std_logic_vector(to_unsigned( 66, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 220, 8)),
16 => std_logic_vector(to_unsigned( 243, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 45, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 687 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 96, 8)),
3 => std_logic_vector(to_unsigned( 241, 8)),
4 => std_logic_vector(to_unsigned( 126, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 225, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 31, 8)),
12 => std_logic_vector(to_unsigned( 119, 8)),
13 => std_logic_vector(to_unsigned( 69, 8)),
14 => std_logic_vector(to_unsigned( 195, 8)),
15 => std_logic_vector(to_unsigned( 84, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110000
elsif count = 688 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 176, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 173, 8)),
5 => std_logic_vector(to_unsigned( 43, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 15, 8)),
10 => std_logic_vector(to_unsigned( 137, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 204, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 221, 8)),
15 => std_logic_vector(to_unsigned( 148, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 204, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 689 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 205, 8)),
3 => std_logic_vector(to_unsigned( 63, 8)),
4 => std_logic_vector(to_unsigned( 30, 8)),
5 => std_logic_vector(to_unsigned( 186, 8)),
6 => std_logic_vector(to_unsigned( 127, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 107, 8)),
10 => std_logic_vector(to_unsigned( 142, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 213, 8)),
13 => std_logic_vector(to_unsigned( 189, 8)),
14 => std_logic_vector(to_unsigned( 174, 8)),
15 => std_logic_vector(to_unsigned( 244, 8)),
16 => std_logic_vector(to_unsigned( 59, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 690 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 37, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 235, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 29, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 156, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 97, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 691 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 234, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 252, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 87, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 132, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 80, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 108, 8)),
16 => std_logic_vector(to_unsigned( 193, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101010
elsif count = 692 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 11, 8)),
3 => std_logic_vector(to_unsigned( 33, 8)),
4 => std_logic_vector(to_unsigned( 205, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 26, 8)),
13 => std_logic_vector(to_unsigned( 45, 8)),
14 => std_logic_vector(to_unsigned( 212, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101101
elsif count = 693 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 22, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 175, 8)),
11 => std_logic_vector(to_unsigned( 225, 8)),
12 => std_logic_vector(to_unsigned( 98, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 7, 8)),
16 => std_logic_vector(to_unsigned( 199, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 694 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 191, 8)),
3 => std_logic_vector(to_unsigned( 232, 8)),
4 => std_logic_vector(to_unsigned( 199, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 45, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 66, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 163, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 125, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 695 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 180, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 189, 8)),
13 => std_logic_vector(to_unsigned( 246, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 89, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 696 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 144, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 66, 8)),
6 => std_logic_vector(to_unsigned( 199, 8)),
7 => std_logic_vector(to_unsigned( 170, 8)),
8 => std_logic_vector(to_unsigned( 15, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 225, 8)),
13 => std_logic_vector(to_unsigned( 48, 8)),
14 => std_logic_vector(to_unsigned( 245, 8)),
15 => std_logic_vector(to_unsigned( 91, 8)),
16 => std_logic_vector(to_unsigned( 254, 8)),
17 => std_logic_vector(to_unsigned( 48, 8)),
18 => std_logic_vector(to_unsigned( 213, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 697 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 116, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 159, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 12, 8)),
9 => std_logic_vector(to_unsigned( 96, 8)),
10 => std_logic_vector(to_unsigned( 188, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 173, 8)),
13 => std_logic_vector(to_unsigned( 176, 8)),
14 => std_logic_vector(to_unsigned( 175, 8)),
15 => std_logic_vector(to_unsigned( 244, 8)),
16 => std_logic_vector(to_unsigned( 58, 8)),
17 => std_logic_vector(to_unsigned( 123, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110011
elsif count = 698 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 51, 8)),
3 => std_logic_vector(to_unsigned( 226, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 117, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 59, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 33, 8)),
12 => std_logic_vector(to_unsigned( 119, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 80, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 179, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 699 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 31, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 77, 8)),
8 => std_logic_vector(to_unsigned( 4, 8)),
9 => std_logic_vector(to_unsigned( 111, 8)),
10 => std_logic_vector(to_unsigned( 104, 8)),
11 => std_logic_vector(to_unsigned( 43, 8)),
12 => std_logic_vector(to_unsigned( 124, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 236, 8)),
17 => std_logic_vector(to_unsigned( 94, 8)),
18 => std_logic_vector(to_unsigned( 162, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010100
elsif count = 700 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 85, 8)),
2 => std_logic_vector(to_unsigned( 157, 8)),
3 => std_logic_vector(to_unsigned( 205, 8)),
4 => std_logic_vector(to_unsigned( 95, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 10, 8)),
8 => std_logic_vector(to_unsigned( 85, 8)),
9 => std_logic_vector(to_unsigned( 97, 8)),
10 => std_logic_vector(to_unsigned( 247, 8)),
11 => std_logic_vector(to_unsigned( 78, 8)),
12 => std_logic_vector(to_unsigned( 246, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 234, 8)),
15 => std_logic_vector(to_unsigned( 107, 8)),
16 => std_logic_vector(to_unsigned( 143, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 701 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 109, 8)),
3 => std_logic_vector(to_unsigned( 242, 8)),
4 => std_logic_vector(to_unsigned( 85, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 206, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 179, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 212, 8)),
13 => std_logic_vector(to_unsigned( 197, 8)),
14 => std_logic_vector(to_unsigned( 141, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 45, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011101
elsif count = 702 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 130, 8)),
2 => std_logic_vector(to_unsigned( 105, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 152, 8)),
6 => std_logic_vector(to_unsigned( 127, 8)),
7 => std_logic_vector(to_unsigned( 171, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 44, 8)),
11 => std_logic_vector(to_unsigned( 94, 8)),
12 => std_logic_vector(to_unsigned( 25, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 48, 8)),
17 => std_logic_vector(to_unsigned( 187, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 703 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 234, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 181, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 48, 8)),
6 => std_logic_vector(to_unsigned( 79, 8)),
7 => std_logic_vector(to_unsigned( 42, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 64, 8)),
11 => std_logic_vector(to_unsigned( 168, 8)),
12 => std_logic_vector(to_unsigned( 71, 8)),
13 => std_logic_vector(to_unsigned( 200, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 25, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 704 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 121, 8)),
3 => std_logic_vector(to_unsigned( 213, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 96, 8)),
10 => std_logic_vector(to_unsigned( 117, 8)),
11 => std_logic_vector(to_unsigned( 201, 8)),
12 => std_logic_vector(to_unsigned( 80, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 68, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 705 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 141, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 128, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 225, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 224, 8)),
13 => std_logic_vector(to_unsigned( 185, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 197, 8)),
16 => std_logic_vector(to_unsigned( 20, 8)),
17 => std_logic_vector(to_unsigned( 73, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 706 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 174, 8)),
2 => std_logic_vector(to_unsigned( 225, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 195, 8)),
5 => std_logic_vector(to_unsigned( 212, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 162, 8)),
11 => std_logic_vector(to_unsigned( 176, 8)),
12 => std_logic_vector(to_unsigned( 76, 8)),
13 => std_logic_vector(to_unsigned( 22, 8)),
14 => std_logic_vector(to_unsigned( 189, 8)),
15 => std_logic_vector(to_unsigned( 8, 8)),
16 => std_logic_vector(to_unsigned( 32, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 186, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 707 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 153, 8)),
7 => std_logic_vector(to_unsigned( 216, 8)),
8 => std_logic_vector(to_unsigned( 53, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 77, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 5, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 180, 8)),
16 => std_logic_vector(to_unsigned( 222, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 82, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 708 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 180, 8)),
2 => std_logic_vector(to_unsigned( 181, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 140, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 117, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 91, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 213, 8)),
12 => std_logic_vector(to_unsigned( 160, 8)),
13 => std_logic_vector(to_unsigned( 211, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 37, 8)),
16 => std_logic_vector(to_unsigned( 225, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 139, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101111
elsif count = 709 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 230, 8)),
2 => std_logic_vector(to_unsigned( 214, 8)),
3 => std_logic_vector(to_unsigned( 89, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 10, 8)),
6 => std_logic_vector(to_unsigned( 14, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 165, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 160, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 215, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 126, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 710 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 228, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 52, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 222, 8)),
8 => std_logic_vector(to_unsigned( 97, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 90, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 47, 8)),
15 => std_logic_vector(to_unsigned( 103, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 711 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 9, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 17, 8)),
4 => std_logic_vector(to_unsigned( 164, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 201, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 137, 8)),
10 => std_logic_vector(to_unsigned( 190, 8)),
11 => std_logic_vector(to_unsigned( 3, 8)),
12 => std_logic_vector(to_unsigned( 182, 8)),
13 => std_logic_vector(to_unsigned( 243, 8)),
14 => std_logic_vector(to_unsigned( 19, 8)),
15 => std_logic_vector(to_unsigned( 44, 8)),
16 => std_logic_vector(to_unsigned( 31, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 180, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 712 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 211, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 240, 8)),
9 => std_logic_vector(to_unsigned( 228, 8)),
10 => std_logic_vector(to_unsigned( 197, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 198, 8)),
13 => std_logic_vector(to_unsigned( 156, 8)),
14 => std_logic_vector(to_unsigned( 185, 8)),
15 => std_logic_vector(to_unsigned( 250, 8)),
16 => std_logic_vector(to_unsigned( 216, 8)),
17 => std_logic_vector(to_unsigned( 192, 8)),
18 => std_logic_vector(to_unsigned( 191, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 713 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 69, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 80, 8)),
5 => std_logic_vector(to_unsigned( 109, 8)),
6 => std_logic_vector(to_unsigned( 31, 8)),
7 => std_logic_vector(to_unsigned( 37, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 48, 8)),
11 => std_logic_vector(to_unsigned( 240, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 136, 8)),
16 => std_logic_vector(to_unsigned( 8, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 43, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 714 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 83, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 185, 8)),
10 => std_logic_vector(to_unsigned( 224, 8)),
11 => std_logic_vector(to_unsigned( 227, 8)),
12 => std_logic_vector(to_unsigned( 182, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 118, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 715 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 48, 8)),
2 => std_logic_vector(to_unsigned( 179, 8)),
3 => std_logic_vector(to_unsigned( 47, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 161, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 111, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 181, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 152, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 207, 8)),
16 => std_logic_vector(to_unsigned( 153, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 716 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 185, 8)),
3 => std_logic_vector(to_unsigned( 7, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 175, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 82, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 78, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 244, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 717 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 27, 8)),
3 => std_logic_vector(to_unsigned( 222, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 158, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 137, 8)),
10 => std_logic_vector(to_unsigned( 77, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 143, 8)),
16 => std_logic_vector(to_unsigned( 71, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 718 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 35, 8)),
2 => std_logic_vector(to_unsigned( 25, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 242, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 212, 8)),
8 => std_logic_vector(to_unsigned( 21, 8)),
9 => std_logic_vector(to_unsigned( 228, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 231, 8)),
12 => std_logic_vector(to_unsigned( 40, 8)),
13 => std_logic_vector(to_unsigned( 185, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 51, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 719 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 68, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 227, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 197, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 220, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 58, 8)),
13 => std_logic_vector(to_unsigned( 49, 8)),
14 => std_logic_vector(to_unsigned( 91, 8)),
15 => std_logic_vector(to_unsigned( 191, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 197, 8)),
18 => std_logic_vector(to_unsigned( 52, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 720 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 101, 8)),
2 => std_logic_vector(to_unsigned( 242, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 72, 8)),
5 => std_logic_vector(to_unsigned( 102, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 89, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 20, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 48, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 721 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 42, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 68, 8)),
4 => std_logic_vector(to_unsigned( 78, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 137, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 249, 8)),
10 => std_logic_vector(to_unsigned( 116, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 119, 8)),
13 => std_logic_vector(to_unsigned( 51, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 121, 8)),
17 => std_logic_vector(to_unsigned( 76, 8)),
18 => std_logic_vector(to_unsigned( 106, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 722 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 94, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 76, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 57, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 13, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 71, 8)),
12 => std_logic_vector(to_unsigned( 179, 8)),
13 => std_logic_vector(to_unsigned( 5, 8)),
14 => std_logic_vector(to_unsigned( 202, 8)),
15 => std_logic_vector(to_unsigned( 25, 8)),
16 => std_logic_vector(to_unsigned( 145, 8)),
17 => std_logic_vector(to_unsigned( 42, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 723 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 163, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 155, 8)),
4 => std_logic_vector(to_unsigned( 47, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 47, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 40, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 38, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 64, 8)),
13 => std_logic_vector(to_unsigned( 38, 8)),
14 => std_logic_vector(to_unsigned( 16, 8)),
15 => std_logic_vector(to_unsigned( 8, 8)),
16 => std_logic_vector(to_unsigned( 20, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 724 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 224, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 153, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 46, 8)),
7 => std_logic_vector(to_unsigned( 189, 8)),
8 => std_logic_vector(to_unsigned( 0, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 153, 8)),
12 => std_logic_vector(to_unsigned( 172, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 66, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 725 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 179, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 14, 8)),
4 => std_logic_vector(to_unsigned( 64, 8)),
5 => std_logic_vector(to_unsigned( 207, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 51, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 67, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 206, 8)),
12 => std_logic_vector(to_unsigned( 108, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 726 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 28, 8)),
4 => std_logic_vector(to_unsigned( 200, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 251, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 198, 8)),
9 => std_logic_vector(to_unsigned( 56, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 105, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 157, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 58, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 727 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 230, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 107, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 4, 8)),
7 => std_logic_vector(to_unsigned( 33, 8)),
8 => std_logic_vector(to_unsigned( 165, 8)),
9 => std_logic_vector(to_unsigned( 222, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 221, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 146, 8)),
15 => std_logic_vector(to_unsigned( 150, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010011
elsif count = 728 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 178, 8)),
5 => std_logic_vector(to_unsigned( 235, 8)),
6 => std_logic_vector(to_unsigned( 190, 8)),
7 => std_logic_vector(to_unsigned( 132, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 180, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 176, 8)),
13 => std_logic_vector(to_unsigned( 95, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 86, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 145, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011000
elsif count = 729 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 25, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 4, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 37, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 64, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 83, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 58, 8)),
14 => std_logic_vector(to_unsigned( 0, 8)),
15 => std_logic_vector(to_unsigned( 35, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 35, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 730 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 119, 8)),
2 => std_logic_vector(to_unsigned( 153, 8)),
3 => std_logic_vector(to_unsigned( 140, 8)),
4 => std_logic_vector(to_unsigned( 174, 8)),
5 => std_logic_vector(to_unsigned( 52, 8)),
6 => std_logic_vector(to_unsigned( 2, 8)),
7 => std_logic_vector(to_unsigned( 87, 8)),
8 => std_logic_vector(to_unsigned( 217, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 156, 8)),
11 => std_logic_vector(to_unsigned( 149, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 108, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 156, 8)),
17 => std_logic_vector(to_unsigned( 142, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 731 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 207, 8)),
2 => std_logic_vector(to_unsigned( 143, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 158, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 182, 8)),
13 => std_logic_vector(to_unsigned( 190, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 93, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 164, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 732 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 219, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 171, 8)),
5 => std_logic_vector(to_unsigned( 117, 8)),
6 => std_logic_vector(to_unsigned( 208, 8)),
7 => std_logic_vector(to_unsigned( 207, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 136, 8)),
10 => std_logic_vector(to_unsigned( 47, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 168, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 221, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 733 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 65, 8)),
7 => std_logic_vector(to_unsigned( 232, 8)),
8 => std_logic_vector(to_unsigned( 241, 8)),
9 => std_logic_vector(to_unsigned( 219, 8)),
10 => std_logic_vector(to_unsigned( 28, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 734 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 235, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 81, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 33, 8)),
7 => std_logic_vector(to_unsigned( 191, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 164, 8)),
11 => std_logic_vector(to_unsigned( 10, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 214, 8)),
15 => std_logic_vector(to_unsigned( 183, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001110
elsif count = 735 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 74, 8)),
2 => std_logic_vector(to_unsigned( 152, 8)),
3 => std_logic_vector(to_unsigned( 166, 8)),
4 => std_logic_vector(to_unsigned( 57, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 78, 8)),
7 => std_logic_vector(to_unsigned( 128, 8)),
8 => std_logic_vector(to_unsigned( 200, 8)),
9 => std_logic_vector(to_unsigned( 200, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 220, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 19, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 736 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 133, 8)),
3 => std_logic_vector(to_unsigned( 244, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 131, 8)),
6 => std_logic_vector(to_unsigned( 66, 8)),
7 => std_logic_vector(to_unsigned( 8, 8)),
8 => std_logic_vector(to_unsigned( 31, 8)),
9 => std_logic_vector(to_unsigned( 101, 8)),
10 => std_logic_vector(to_unsigned( 168, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 189, 8)),
13 => std_logic_vector(to_unsigned( 239, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 162, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 737 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 87, 8)),
7 => std_logic_vector(to_unsigned( 180, 8)),
8 => std_logic_vector(to_unsigned( 169, 8)),
9 => std_logic_vector(to_unsigned( 143, 8)),
10 => std_logic_vector(to_unsigned( 200, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 36, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 49, 8)),
16 => std_logic_vector(to_unsigned( 240, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 738 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 195, 8)),
2 => std_logic_vector(to_unsigned( 91, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 232, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 61, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 225, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 28, 8)),
11 => std_logic_vector(to_unsigned( 55, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 187, 8)),
16 => std_logic_vector(to_unsigned( 83, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 739 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 38, 8)),
3 => std_logic_vector(to_unsigned( 133, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 133, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 229, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 26, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 157, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 197, 8)),
16 => std_logic_vector(to_unsigned( 206, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 740 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 226, 8)),
3 => std_logic_vector(to_unsigned( 209, 8)),
4 => std_logic_vector(to_unsigned( 184, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 36, 8)),
7 => std_logic_vector(to_unsigned( 31, 8)),
8 => std_logic_vector(to_unsigned( 103, 8)),
9 => std_logic_vector(to_unsigned( 35, 8)),
10 => std_logic_vector(to_unsigned( 63, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 53, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 36, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 741 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 253, 8)),
2 => std_logic_vector(to_unsigned( 13, 8)),
3 => std_logic_vector(to_unsigned( 154, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 131, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 95, 8)),
11 => std_logic_vector(to_unsigned( 46, 8)),
12 => std_logic_vector(to_unsigned( 50, 8)),
13 => std_logic_vector(to_unsigned( 160, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 231, 8)),
16 => std_logic_vector(to_unsigned( 5, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 742 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 57, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 21, 8)),
4 => std_logic_vector(to_unsigned( 47, 8)),
5 => std_logic_vector(to_unsigned( 27, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 77, 8)),
9 => std_logic_vector(to_unsigned( 224, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 92, 8)),
12 => std_logic_vector(to_unsigned( 48, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 33, 8)),
15 => std_logic_vector(to_unsigned( 45, 8)),
16 => std_logic_vector(to_unsigned( 37, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 743 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 158, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 245, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 211, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 83, 8)),
17 => std_logic_vector(to_unsigned( 196, 8)),
18 => std_logic_vector(to_unsigned( 119, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101001
elsif count = 744 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 34, 8)),
3 => std_logic_vector(to_unsigned( 128, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 117, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 187, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 27, 8)),
11 => std_logic_vector(to_unsigned( 76, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 77, 8)),
16 => std_logic_vector(to_unsigned( 157, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 745 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 216, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 38, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 84, 8)),
7 => std_logic_vector(to_unsigned( 77, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 53, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 127, 8)),
12 => std_logic_vector(to_unsigned( 192, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 56, 8)),
15 => std_logic_vector(to_unsigned( 178, 8)),
16 => std_logic_vector(to_unsigned( 60, 8)),
17 => std_logic_vector(to_unsigned( 108, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111100
elsif count = 746 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 195, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 238, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 136, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 78, 8)),
11 => std_logic_vector(to_unsigned( 125, 8)),
12 => std_logic_vector(to_unsigned( 228, 8)),
13 => std_logic_vector(to_unsigned( 246, 8)),
14 => std_logic_vector(to_unsigned( 8, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 244, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 747 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 166, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 195, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 230, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 179, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 175, 8)),
13 => std_logic_vector(to_unsigned( 202, 8)),
14 => std_logic_vector(to_unsigned( 51, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 748 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 6, 8)),
2 => std_logic_vector(to_unsigned( 15, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 7, 8)),
5 => std_logic_vector(to_unsigned( 123, 8)),
6 => std_logic_vector(to_unsigned( 44, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 202, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 58, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 131, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 237, 8)),
17 => std_logic_vector(to_unsigned( 151, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011000
elsif count = 749 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 16, 8)),
2 => std_logic_vector(to_unsigned( 0, 8)),
3 => std_logic_vector(to_unsigned( 200, 8)),
4 => std_logic_vector(to_unsigned( 221, 8)),
5 => std_logic_vector(to_unsigned( 248, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 215, 8)),
8 => std_logic_vector(to_unsigned( 206, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 160, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 27, 8)),
14 => std_logic_vector(to_unsigned( 22, 8)),
15 => std_logic_vector(to_unsigned( 198, 8)),
16 => std_logic_vector(to_unsigned( 223, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 750 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 45, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 177, 8)),
5 => std_logic_vector(to_unsigned( 232, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 139, 8)),
10 => std_logic_vector(to_unsigned( 224, 8)),
11 => std_logic_vector(to_unsigned( 53, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 208, 8)),
15 => std_logic_vector(to_unsigned( 50, 8)),
16 => std_logic_vector(to_unsigned( 34, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 751 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 59, 8)),
2 => std_logic_vector(to_unsigned( 1, 8)),
3 => std_logic_vector(to_unsigned( 37, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 32, 8)),
7 => std_logic_vector(to_unsigned( 254, 8)),
8 => std_logic_vector(to_unsigned( 228, 8)),
9 => std_logic_vector(to_unsigned( 145, 8)),
10 => std_logic_vector(to_unsigned( 87, 8)),
11 => std_logic_vector(to_unsigned( 14, 8)),
12 => std_logic_vector(to_unsigned( 104, 8)),
13 => std_logic_vector(to_unsigned( 159, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110010
elsif count = 752 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 176, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 238, 8)),
5 => std_logic_vector(to_unsigned( 118, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 165, 8)),
9 => std_logic_vector(to_unsigned( 145, 8)),
10 => std_logic_vector(to_unsigned( 214, 8)),
11 => std_logic_vector(to_unsigned( 106, 8)),
12 => std_logic_vector(to_unsigned( 227, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 202, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 753 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 111, 8)),
4 => std_logic_vector(to_unsigned( 229, 8)),
5 => std_logic_vector(to_unsigned( 43, 8)),
6 => std_logic_vector(to_unsigned( 156, 8)),
7 => std_logic_vector(to_unsigned( 160, 8)),
8 => std_logic_vector(to_unsigned( 231, 8)),
9 => std_logic_vector(to_unsigned( 148, 8)),
10 => std_logic_vector(to_unsigned( 111, 8)),
11 => std_logic_vector(to_unsigned( 34, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 60, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 754 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 16, 8)),
2 => std_logic_vector(to_unsigned( 128, 8)),
3 => std_logic_vector(to_unsigned( 166, 8)),
4 => std_logic_vector(to_unsigned( 192, 8)),
5 => std_logic_vector(to_unsigned( 99, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 69, 8)),
9 => std_logic_vector(to_unsigned( 188, 8)),
10 => std_logic_vector(to_unsigned( 18, 8)),
11 => std_logic_vector(to_unsigned( 8, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 9, 8)),
17 => std_logic_vector(to_unsigned( 79, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 755 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 66, 8)),
2 => std_logic_vector(to_unsigned( 93, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 89, 8)),
7 => std_logic_vector(to_unsigned( 38, 8)),
8 => std_logic_vector(to_unsigned( 48, 8)),
9 => std_logic_vector(to_unsigned( 208, 8)),
10 => std_logic_vector(to_unsigned( 239, 8)),
11 => std_logic_vector(to_unsigned( 95, 8)),
12 => std_logic_vector(to_unsigned( 214, 8)),
13 => std_logic_vector(to_unsigned( 78, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 104, 8)),
16 => std_logic_vector(to_unsigned( 205, 8)),
17 => std_logic_vector(to_unsigned( 78, 8)),
18 => std_logic_vector(to_unsigned( 156, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 756 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 116, 8)),
2 => std_logic_vector(to_unsigned( 198, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 209, 8)),
6 => std_logic_vector(to_unsigned( 126, 8)),
7 => std_logic_vector(to_unsigned( 16, 8)),
8 => std_logic_vector(to_unsigned( 205, 8)),
9 => std_logic_vector(to_unsigned( 188, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 219, 8)),
12 => std_logic_vector(to_unsigned( 23, 8)),
13 => std_logic_vector(to_unsigned( 151, 8)),
14 => std_logic_vector(to_unsigned( 116, 8)),
15 => std_logic_vector(to_unsigned( 157, 8)),
16 => std_logic_vector(to_unsigned( 108, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 115, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 757 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 175, 8)),
3 => std_logic_vector(to_unsigned( 239, 8)),
4 => std_logic_vector(to_unsigned( 106, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 66, 8)),
7 => std_logic_vector(to_unsigned( 178, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 219, 8)),
10 => std_logic_vector(to_unsigned( 126, 8)),
11 => std_logic_vector(to_unsigned( 1, 8)),
12 => std_logic_vector(to_unsigned( 95, 8)),
13 => std_logic_vector(to_unsigned( 209, 8)),
14 => std_logic_vector(to_unsigned( 62, 8)),
15 => std_logic_vector(to_unsigned( 4, 8)),
16 => std_logic_vector(to_unsigned( 186, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 758 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 139, 8)),
2 => std_logic_vector(to_unsigned( 23, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 234, 8)),
5 => std_logic_vector(to_unsigned( 129, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 38, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 35, 8)),
12 => std_logic_vector(to_unsigned( 160, 8)),
13 => std_logic_vector(to_unsigned( 51, 8)),
14 => std_logic_vector(to_unsigned( 208, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 215, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110000
elsif count = 759 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 74, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 180, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 16, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 206, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 147, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 760 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 165, 8)),
3 => std_logic_vector(to_unsigned( 12, 8)),
4 => std_logic_vector(to_unsigned( 39, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 9, 8)),
7 => std_logic_vector(to_unsigned( 11, 8)),
8 => std_logic_vector(to_unsigned( 7, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 168, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 251, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 229, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110001
elsif count = 761 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 136, 8)),
4 => std_logic_vector(to_unsigned( 52, 8)),
5 => std_logic_vector(to_unsigned( 120, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 139, 8)),
8 => std_logic_vector(to_unsigned( 33, 8)),
9 => std_logic_vector(to_unsigned( 114, 8)),
10 => std_logic_vector(to_unsigned( 70, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 167, 8)),
14 => std_logic_vector(to_unsigned( 216, 8)),
15 => std_logic_vector(to_unsigned( 123, 8)),
16 => std_logic_vector(to_unsigned( 61, 8)),
17 => std_logic_vector(to_unsigned( 134, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 762 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 224, 8)),
6 => std_logic_vector(to_unsigned( 241, 8)),
7 => std_logic_vector(to_unsigned( 128, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 167, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 154, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 189, 8)),
15 => std_logic_vector(to_unsigned( 39, 8)),
16 => std_logic_vector(to_unsigned( 84, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111010
elsif count = 763 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 41, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 74, 8)),
4 => std_logic_vector(to_unsigned( 43, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 76, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 61, 8)),
10 => std_logic_vector(to_unsigned( 48, 8)),
11 => std_logic_vector(to_unsigned( 251, 8)),
12 => std_logic_vector(to_unsigned( 90, 8)),
13 => std_logic_vector(to_unsigned( 33, 8)),
14 => std_logic_vector(to_unsigned( 94, 8)),
15 => std_logic_vector(to_unsigned( 45, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 764 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 198, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 181, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 159, 8)),
8 => std_logic_vector(to_unsigned( 197, 8)),
9 => std_logic_vector(to_unsigned( 85, 8)),
10 => std_logic_vector(to_unsigned( 123, 8)),
11 => std_logic_vector(to_unsigned( 211, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 42, 8)),
16 => std_logic_vector(to_unsigned( 231, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 765 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 103, 8)),
2 => std_logic_vector(to_unsigned( 145, 8)),
3 => std_logic_vector(to_unsigned( 19, 8)),
4 => std_logic_vector(to_unsigned( 33, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 225, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 148, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 214, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 227, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 193, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 766 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 42, 8)),
2 => std_logic_vector(to_unsigned( 67, 8)),
3 => std_logic_vector(to_unsigned( 191, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 70, 8)),
7 => std_logic_vector(to_unsigned( 254, 8)),
8 => std_logic_vector(to_unsigned( 54, 8)),
9 => std_logic_vector(to_unsigned( 78, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 42, 8)),
13 => std_logic_vector(to_unsigned( 77, 8)),
14 => std_logic_vector(to_unsigned( 42, 8)),
15 => std_logic_vector(to_unsigned( 241, 8)),
16 => std_logic_vector(to_unsigned( 252, 8)),
17 => std_logic_vector(to_unsigned( 47, 8)),
18 => std_logic_vector(to_unsigned( 36, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 767 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 113, 8)),
2 => std_logic_vector(to_unsigned( 25, 8)),
3 => std_logic_vector(to_unsigned( 85, 8)),
4 => std_logic_vector(to_unsigned( 29, 8)),
5 => std_logic_vector(to_unsigned( 137, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 34, 8)),
9 => std_logic_vector(to_unsigned( 223, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 66, 8)),
12 => std_logic_vector(to_unsigned( 52, 8)),
13 => std_logic_vector(to_unsigned( 201, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 79, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 50, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 768 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 113, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 13, 8)),
9 => std_logic_vector(to_unsigned( 251, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 114, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 769 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 56, 8)),
2 => std_logic_vector(to_unsigned( 117, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 53, 8)),
5 => std_logic_vector(to_unsigned( 100, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 88, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 86, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 166, 8)),
14 => std_logic_vector(to_unsigned( 64, 8)),
15 => std_logic_vector(to_unsigned( 208, 8)),
16 => std_logic_vector(to_unsigned( 239, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 770 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 121, 8)),
3 => std_logic_vector(to_unsigned( 4, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 156, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 80, 8)),
9 => std_logic_vector(to_unsigned( 199, 8)),
10 => std_logic_vector(to_unsigned( 245, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 138, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 146, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 771 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 50, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 86, 8)),
4 => std_logic_vector(to_unsigned( 132, 8)),
5 => std_logic_vector(to_unsigned( 40, 8)),
6 => std_logic_vector(to_unsigned( 174, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 171, 8)),
9 => std_logic_vector(to_unsigned( 59, 8)),
10 => std_logic_vector(to_unsigned( 117, 8)),
11 => std_logic_vector(to_unsigned( 37, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 58, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 231, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 772 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 134, 8)),
3 => std_logic_vector(to_unsigned( 143, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 59, 8)),
6 => std_logic_vector(to_unsigned( 127, 8)),
7 => std_logic_vector(to_unsigned( 53, 8)),
8 => std_logic_vector(to_unsigned( 59, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 55, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 57, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 773 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 117, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 203, 8)),
4 => std_logic_vector(to_unsigned( 73, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 112, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 104, 8)),
10 => std_logic_vector(to_unsigned( 89, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 79, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 35, 8)),
15 => std_logic_vector(to_unsigned( 15, 8)),
16 => std_logic_vector(to_unsigned( 197, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 62, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110001
elsif count = 774 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 92, 8)),
2 => std_logic_vector(to_unsigned( 80, 8)),
3 => std_logic_vector(to_unsigned( 134, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 18, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 21, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 143, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 141, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 96, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 775 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 247, 8)),
4 => std_logic_vector(to_unsigned( 92, 8)),
5 => std_logic_vector(to_unsigned( 43, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 56, 8)),
8 => std_logic_vector(to_unsigned( 191, 8)),
9 => std_logic_vector(to_unsigned( 94, 8)),
10 => std_logic_vector(to_unsigned( 173, 8)),
11 => std_logic_vector(to_unsigned( 176, 8)),
12 => std_logic_vector(to_unsigned( 66, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 87, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 170, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 776 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 14, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 156, 8)),
4 => std_logic_vector(to_unsigned( 197, 8)),
5 => std_logic_vector(to_unsigned( 103, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 239, 8)),
12 => std_logic_vector(to_unsigned( 42, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 169, 8)),
16 => std_logic_vector(to_unsigned( 128, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 777 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 120, 8)),
2 => std_logic_vector(to_unsigned( 201, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 203, 8)),
5 => std_logic_vector(to_unsigned( 229, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 115, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 238, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 16, 8)),
16 => std_logic_vector(to_unsigned( 47, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 778 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 209, 8)),
2 => std_logic_vector(to_unsigned( 31, 8)),
3 => std_logic_vector(to_unsigned( 184, 8)),
4 => std_logic_vector(to_unsigned( 130, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 159, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 95, 8)),
12 => std_logic_vector(to_unsigned( 129, 8)),
13 => std_logic_vector(to_unsigned( 228, 8)),
14 => std_logic_vector(to_unsigned( 242, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 139, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 779 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 186, 8)),
2 => std_logic_vector(to_unsigned( 67, 8)),
3 => std_logic_vector(to_unsigned( 226, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 184, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 202, 8)),
8 => std_logic_vector(to_unsigned( 123, 8)),
9 => std_logic_vector(to_unsigned( 167, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 186, 8)),
12 => std_logic_vector(to_unsigned( 67, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 212, 8)),
15 => std_logic_vector(to_unsigned( 188, 8)),
16 => std_logic_vector(to_unsigned( 65, 8)),
17 => std_logic_vector(to_unsigned( 197, 8)),
18 => std_logic_vector(to_unsigned( 92, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111101
elsif count = 780 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 168, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 215, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 22, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 24, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 57, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 153, 8)),
15 => std_logic_vector(to_unsigned( 56, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101000
elsif count = 781 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 142, 8)),
3 => std_logic_vector(to_unsigned( 229, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 20, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 101, 8)),
17 => std_logic_vector(to_unsigned( 130, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011001
elsif count = 782 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 249, 8)),
2 => std_logic_vector(to_unsigned( 35, 8)),
3 => std_logic_vector(to_unsigned( 174, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 167, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 69, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 106, 8)),
11 => std_logic_vector(to_unsigned( 98, 8)),
12 => std_logic_vector(to_unsigned( 110, 8)),
13 => std_logic_vector(to_unsigned( 127, 8)),
14 => std_logic_vector(to_unsigned( 16, 8)),
15 => std_logic_vector(to_unsigned( 64, 8)),
16 => std_logic_vector(to_unsigned( 28, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111000
elsif count = 783 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 33, 8)),
2 => std_logic_vector(to_unsigned( 52, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 53, 8)),
5 => std_logic_vector(to_unsigned( 191, 8)),
6 => std_logic_vector(to_unsigned( 239, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 43, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 38, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 21, 8)),
15 => std_logic_vector(to_unsigned( 54, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 78, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111011
elsif count = 784 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 137, 8)),
3 => std_logic_vector(to_unsigned( 145, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 229, 8)),
6 => std_logic_vector(to_unsigned( 101, 8)),
7 => std_logic_vector(to_unsigned( 199, 8)),
8 => std_logic_vector(to_unsigned( 137, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 75, 8)),
11 => std_logic_vector(to_unsigned( 153, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 176, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 36, 8)),
16 => std_logic_vector(to_unsigned( 15, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 785 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 122, 8)),
2 => std_logic_vector(to_unsigned( 204, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 142, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 106, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 209, 8)),
11 => std_logic_vector(to_unsigned( 123, 8)),
12 => std_logic_vector(to_unsigned( 158, 8)),
13 => std_logic_vector(to_unsigned( 2, 8)),
14 => std_logic_vector(to_unsigned( 193, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111110
elsif count = 786 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 133, 8)),
2 => std_logic_vector(to_unsigned( 47, 8)),
3 => std_logic_vector(to_unsigned( 151, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 203, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 20, 8)),
8 => std_logic_vector(to_unsigned( 4, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 166, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 27, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 787 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 238, 8)),
6 => std_logic_vector(to_unsigned( 104, 8)),
7 => std_logic_vector(to_unsigned( 46, 8)),
8 => std_logic_vector(to_unsigned( 90, 8)),
9 => std_logic_vector(to_unsigned( 183, 8)),
10 => std_logic_vector(to_unsigned( 180, 8)),
11 => std_logic_vector(to_unsigned( 130, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 121, 8)),
14 => std_logic_vector(to_unsigned( 137, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 788 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 29, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 165, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 95, 8)),
6 => std_logic_vector(to_unsigned( 117, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 87, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 158, 8)),
12 => std_logic_vector(to_unsigned( 168, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 179, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 789 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 89, 8)),
2 => std_logic_vector(to_unsigned( 201, 8)),
3 => std_logic_vector(to_unsigned( 246, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 29, 8)),
7 => std_logic_vector(to_unsigned( 78, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 111, 8)),
12 => std_logic_vector(to_unsigned( 17, 8)),
13 => std_logic_vector(to_unsigned( 79, 8)),
14 => std_logic_vector(to_unsigned( 51, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 73, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 42, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 790 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 170, 8)),
3 => std_logic_vector(to_unsigned( 159, 8)),
4 => std_logic_vector(to_unsigned( 158, 8)),
5 => std_logic_vector(to_unsigned( 217, 8)),
6 => std_logic_vector(to_unsigned( 233, 8)),
7 => std_logic_vector(to_unsigned( 34, 8)),
8 => std_logic_vector(to_unsigned( 122, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 23, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 19, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111001
elsif count = 791 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 216, 8)),
3 => std_logic_vector(to_unsigned( 174, 8)),
4 => std_logic_vector(to_unsigned( 216, 8)),
5 => std_logic_vector(to_unsigned( 185, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 198, 8)),
8 => std_logic_vector(to_unsigned( 192, 8)),
9 => std_logic_vector(to_unsigned( 191, 8)),
10 => std_logic_vector(to_unsigned( 85, 8)),
11 => std_logic_vector(to_unsigned( 10, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 195, 8)),
15 => std_logic_vector(to_unsigned( 248, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 792 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 198, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 209, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 210, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 179, 8)),
12 => std_logic_vector(to_unsigned( 240, 8)),
13 => std_logic_vector(to_unsigned( 226, 8)),
14 => std_logic_vector(to_unsigned( 83, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 163, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001110
elsif count = 793 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 58, 8)),
2 => std_logic_vector(to_unsigned( 203, 8)),
3 => std_logic_vector(to_unsigned( 119, 8)),
4 => std_logic_vector(to_unsigned( 222, 8)),
5 => std_logic_vector(to_unsigned( 94, 8)),
6 => std_logic_vector(to_unsigned( 239, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 146, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 189, 8)),
11 => std_logic_vector(to_unsigned( 133, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 224, 8)),
14 => std_logic_vector(to_unsigned( 149, 8)),
15 => std_logic_vector(to_unsigned( 1, 8)),
16 => std_logic_vector(to_unsigned( 78, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 187, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 794 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 230, 8)),
2 => std_logic_vector(to_unsigned( 169, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 33, 8)),
5 => std_logic_vector(to_unsigned( 105, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 181, 8)),
8 => std_logic_vector(to_unsigned( 222, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 114, 8)),
11 => std_logic_vector(to_unsigned( 226, 8)),
12 => std_logic_vector(to_unsigned( 177, 8)),
13 => std_logic_vector(to_unsigned( 153, 8)),
14 => std_logic_vector(to_unsigned( 126, 8)),
15 => std_logic_vector(to_unsigned( 102, 8)),
16 => std_logic_vector(to_unsigned( 22, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 795 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 127, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 195, 8)),
5 => std_logic_vector(to_unsigned( 68, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 3, 8)),
8 => std_logic_vector(to_unsigned( 186, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 103, 8)),
13 => std_logic_vector(to_unsigned( 198, 8)),
14 => std_logic_vector(to_unsigned( 58, 8)),
15 => std_logic_vector(to_unsigned( 25, 8)),
16 => std_logic_vector(to_unsigned( 85, 8)),
17 => std_logic_vector(to_unsigned( 82, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010101
elsif count = 796 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 137, 8)),
8 => std_logic_vector(to_unsigned( 119, 8)),
9 => std_logic_vector(to_unsigned( 124, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 52, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 201, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 797 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 78, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 233, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 55, 8)),
8 => std_logic_vector(to_unsigned( 214, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 94, 8)),
11 => std_logic_vector(to_unsigned( 111, 8)),
12 => std_logic_vector(to_unsigned( 222, 8)),
13 => std_logic_vector(to_unsigned( 5, 8)),
14 => std_logic_vector(to_unsigned( 212, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 203, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 798 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 71, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 142, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 13, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 81, 8)),
10 => std_logic_vector(to_unsigned( 197, 8)),
11 => std_logic_vector(to_unsigned( 67, 8)),
12 => std_logic_vector(to_unsigned( 195, 8)),
13 => std_logic_vector(to_unsigned( 45, 8)),
14 => std_logic_vector(to_unsigned( 205, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 167, 8)),
17 => std_logic_vector(to_unsigned( 75, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 799 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 207, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 167, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 199, 8)),
8 => std_logic_vector(to_unsigned( 191, 8)),
9 => std_logic_vector(to_unsigned( 60, 8)),
10 => std_logic_vector(to_unsigned( 250, 8)),
11 => std_logic_vector(to_unsigned( 28, 8)),
12 => std_logic_vector(to_unsigned( 197, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 213, 8)),
16 => std_logic_vector(to_unsigned( 173, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 175, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 800 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 92, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 40, 8)),
4 => std_logic_vector(to_unsigned( 45, 8)),
5 => std_logic_vector(to_unsigned( 60, 8)),
6 => std_logic_vector(to_unsigned( 25, 8)),
7 => std_logic_vector(to_unsigned( 61, 8)),
8 => std_logic_vector(to_unsigned( 112, 8)),
9 => std_logic_vector(to_unsigned( 98, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 14, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 83, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 2, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011110
elsif count = 801 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 25, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 14, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 249, 8)),
6 => std_logic_vector(to_unsigned( 33, 8)),
7 => std_logic_vector(to_unsigned( 28, 8)),
8 => std_logic_vector(to_unsigned( 175, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 219, 8)),
13 => std_logic_vector(to_unsigned( 52, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001011
elsif count = 802 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 128, 8)),
2 => std_logic_vector(to_unsigned( 72, 8)),
3 => std_logic_vector(to_unsigned( 49, 8)),
4 => std_logic_vector(to_unsigned( 80, 8)),
5 => std_logic_vector(to_unsigned( 89, 8)),
6 => std_logic_vector(to_unsigned( 123, 8)),
7 => std_logic_vector(to_unsigned( 108, 8)),
8 => std_logic_vector(to_unsigned( 60, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 123, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 60, 8)),
15 => std_logic_vector(to_unsigned( 70, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 112, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 803 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 69, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 189, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 156, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 252, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 161, 8)),
15 => std_logic_vector(to_unsigned( 88, 8)),
16 => std_logic_vector(to_unsigned( 77, 8)),
17 => std_logic_vector(to_unsigned( 107, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001101
elsif count = 804 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 202, 8)),
2 => std_logic_vector(to_unsigned( 156, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 163, 8)),
6 => std_logic_vector(to_unsigned( 157, 8)),
7 => std_logic_vector(to_unsigned( 145, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 245, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 140, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 136, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 183, 8)),
18 => std_logic_vector(to_unsigned( 185, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 805 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 242, 8)),
2 => std_logic_vector(to_unsigned( 127, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 158, 8)),
5 => std_logic_vector(to_unsigned( 4, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 139, 8)),
9 => std_logic_vector(to_unsigned( 247, 8)),
10 => std_logic_vector(to_unsigned( 103, 8)),
11 => std_logic_vector(to_unsigned( 137, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 199, 8)),
14 => std_logic_vector(to_unsigned( 165, 8)),
15 => std_logic_vector(to_unsigned( 123, 8)),
16 => std_logic_vector(to_unsigned( 191, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101010
elsif count = 806 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 29, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 216, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 223, 8)),
7 => std_logic_vector(to_unsigned( 253, 8)),
8 => std_logic_vector(to_unsigned( 65, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 98, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 123, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 90, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110101
elsif count = 807 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 181, 8)),
4 => std_logic_vector(to_unsigned( 244, 8)),
5 => std_logic_vector(to_unsigned( 226, 8)),
6 => std_logic_vector(to_unsigned( 23, 8)),
7 => std_logic_vector(to_unsigned( 18, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 231, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 112, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 64, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 199, 8)),
16 => std_logic_vector(to_unsigned( 150, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 188, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 808 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 99, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 123, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 148, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 97, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 47, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 109, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 98, 8)),
15 => std_logic_vector(to_unsigned( 24, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 809 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 173, 8)),
2 => std_logic_vector(to_unsigned( 138, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 107, 8)),
5 => std_logic_vector(to_unsigned( 246, 8)),
6 => std_logic_vector(to_unsigned( 115, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 217, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 28, 8)),
11 => std_logic_vector(to_unsigned( 183, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 12, 8)),
15 => std_logic_vector(to_unsigned( 151, 8)),
16 => std_logic_vector(to_unsigned( 246, 8)),
17 => std_logic_vector(to_unsigned( 117, 8)),
18 => std_logic_vector(to_unsigned( 160, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 810 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 204, 8)),
2 => std_logic_vector(to_unsigned( 200, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 34, 8)),
6 => std_logic_vector(to_unsigned( 9, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 171, 8)),
9 => std_logic_vector(to_unsigned( 47, 8)),
10 => std_logic_vector(to_unsigned( 232, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 208, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 139, 8)),
15 => std_logic_vector(to_unsigned( 16, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 811 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 215, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 36, 8)),
6 => std_logic_vector(to_unsigned( 221, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 214, 8)),
9 => std_logic_vector(to_unsigned( 173, 8)),
10 => std_logic_vector(to_unsigned( 86, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 22, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 154, 8)),
15 => std_logic_vector(to_unsigned( 176, 8)),
16 => std_logic_vector(to_unsigned( 89, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 148, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 812 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 152, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 160, 8)),
4 => std_logic_vector(to_unsigned( 89, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 152, 8)),
7 => std_logic_vector(to_unsigned( 32, 8)),
8 => std_logic_vector(to_unsigned( 73, 8)),
9 => std_logic_vector(to_unsigned( 166, 8)),
10 => std_logic_vector(to_unsigned( 141, 8)),
11 => std_logic_vector(to_unsigned( 68, 8)),
12 => std_logic_vector(to_unsigned( 168, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 19, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 813 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 227, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 57, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 72, 8)),
8 => std_logic_vector(to_unsigned( 209, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 175, 8)),
11 => std_logic_vector(to_unsigned( 217, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 124, 8)),
14 => std_logic_vector(to_unsigned( 213, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 167, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011100
elsif count = 814 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 12, 8)),
2 => std_logic_vector(to_unsigned( 242, 8)),
3 => std_logic_vector(to_unsigned( 50, 8)),
4 => std_logic_vector(to_unsigned( 50, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 44, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 14, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 26, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 66, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 198, 8)),
16 => std_logic_vector(to_unsigned( 50, 8)),
17 => std_logic_vector(to_unsigned( 85, 8)),
18 => std_logic_vector(to_unsigned( 44, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 815 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 26, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 173, 8)),
6 => std_logic_vector(to_unsigned( 161, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 63, 8)),
9 => std_logic_vector(to_unsigned( 170, 8)),
10 => std_logic_vector(to_unsigned( 158, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 172, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 86, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 174, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010110
elsif count = 816 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 196, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 255, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 156, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 214, 8)),
8 => std_logic_vector(to_unsigned( 156, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 162, 8)),
14 => std_logic_vector(to_unsigned( 202, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 24, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 136, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101101
elsif count = 817 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 225, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 105, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 168, 8)),
10 => std_logic_vector(to_unsigned( 215, 8)),
11 => std_logic_vector(to_unsigned( 197, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 236, 8)),
14 => std_logic_vector(to_unsigned( 90, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 202, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 818 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 116, 8)),
2 => std_logic_vector(to_unsigned( 71, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 59, 8)),
5 => std_logic_vector(to_unsigned( 139, 8)),
6 => std_logic_vector(to_unsigned( 94, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 69, 8)),
9 => std_logic_vector(to_unsigned( 62, 8)),
10 => std_logic_vector(to_unsigned( 101, 8)),
11 => std_logic_vector(to_unsigned( 85, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 230, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 127, 8)),
17 => std_logic_vector(to_unsigned( 104, 8)),
18 => std_logic_vector(to_unsigned( 103, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111111
elsif count = 819 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 3, 8)),
2 => std_logic_vector(to_unsigned( 241, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 106, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 80, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 186, 8)),
9 => std_logic_vector(to_unsigned( 121, 8)),
10 => std_logic_vector(to_unsigned( 122, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 140, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 89, 8)),
16 => std_logic_vector(to_unsigned( 68, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110110
elsif count = 820 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 34, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 76, 8)),
4 => std_logic_vector(to_unsigned( 179, 8)),
5 => std_logic_vector(to_unsigned( 42, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 31, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 90, 8)),
12 => std_logic_vector(to_unsigned( 165, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 127, 8)),
16 => std_logic_vector(to_unsigned( 9, 8)),
17 => std_logic_vector(to_unsigned( 57, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 821 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 15, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 20, 8)),
4 => std_logic_vector(to_unsigned( 116, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 77, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 121, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 5, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 111, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 822 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 88, 8)),
2 => std_logic_vector(to_unsigned( 27, 8)),
3 => std_logic_vector(to_unsigned( 131, 8)),
4 => std_logic_vector(to_unsigned( 100, 8)),
5 => std_logic_vector(to_unsigned( 48, 8)),
6 => std_logic_vector(to_unsigned( 45, 8)),
7 => std_logic_vector(to_unsigned( 82, 8)),
8 => std_logic_vector(to_unsigned( 149, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 34, 8)),
12 => std_logic_vector(to_unsigned( 111, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 80, 8)),
16 => std_logic_vector(to_unsigned( 19, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 823 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 202, 8)),
2 => std_logic_vector(to_unsigned( 111, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 214, 8)),
6 => std_logic_vector(to_unsigned( 99, 8)),
7 => std_logic_vector(to_unsigned( 194, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 126, 8)),
10 => std_logic_vector(to_unsigned( 73, 8)),
11 => std_logic_vector(to_unsigned( 135, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 79, 8)),
15 => std_logic_vector(to_unsigned( 136, 8)),
16 => std_logic_vector(to_unsigned( 172, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 824 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 64, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 32, 8)),
8 => std_logic_vector(to_unsigned( 13, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 184, 8)),
12 => std_logic_vector(to_unsigned( 32, 8)),
13 => std_logic_vector(to_unsigned( 200, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 45, 8)),
16 => std_logic_vector(to_unsigned( 125, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110110
elsif count = 825 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 82, 8)),
4 => std_logic_vector(to_unsigned( 150, 8)),
5 => std_logic_vector(to_unsigned( 32, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 8, 8)),
8 => std_logic_vector(to_unsigned( 45, 8)),
9 => std_logic_vector(to_unsigned( 202, 8)),
10 => std_logic_vector(to_unsigned( 10, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 200, 8)),
13 => std_logic_vector(to_unsigned( 58, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 63, 8)),
18 => std_logic_vector(to_unsigned( 122, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 826 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 87, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 182, 8)),
11 => std_logic_vector(to_unsigned( 81, 8)),
12 => std_logic_vector(to_unsigned( 122, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 119, 8)),
15 => std_logic_vector(to_unsigned( 15, 8)),
16 => std_logic_vector(to_unsigned( 177, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 827 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 80, 8)),
2 => std_logic_vector(to_unsigned( 216, 8)),
3 => std_logic_vector(to_unsigned( 66, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 143, 8)),
6 => std_logic_vector(to_unsigned( 187, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 76, 8)),
9 => std_logic_vector(to_unsigned( 161, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 42, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 249, 8)),
16 => std_logic_vector(to_unsigned( 251, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111000
elsif count = 828 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 190, 8)),
5 => std_logic_vector(to_unsigned( 67, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 28, 8)),
8 => std_logic_vector(to_unsigned( 101, 8)),
9 => std_logic_vector(to_unsigned( 92, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 115, 8)),
12 => std_logic_vector(to_unsigned( 14, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 254, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 829 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 186, 8)),
2 => std_logic_vector(to_unsigned( 67, 8)),
3 => std_logic_vector(to_unsigned( 177, 8)),
4 => std_logic_vector(to_unsigned( 175, 8)),
5 => std_logic_vector(to_unsigned( 49, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 145, 8)),
11 => std_logic_vector(to_unsigned( 50, 8)),
12 => std_logic_vector(to_unsigned( 3, 8)),
13 => std_logic_vector(to_unsigned( 218, 8)),
14 => std_logic_vector(to_unsigned( 144, 8)),
15 => std_logic_vector(to_unsigned( 113, 8)),
16 => std_logic_vector(to_unsigned( 177, 8)),
17 => std_logic_vector(to_unsigned( 203, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011010
elsif count = 830 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 178, 8)),
2 => std_logic_vector(to_unsigned( 228, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 203, 8)),
5 => std_logic_vector(to_unsigned( 218, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 175, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 33, 8)),
10 => std_logic_vector(to_unsigned( 171, 8)),
11 => std_logic_vector(to_unsigned( 131, 8)),
12 => std_logic_vector(to_unsigned( 211, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 136, 8)),
17 => std_logic_vector(to_unsigned( 159, 8)),
18 => std_logic_vector(to_unsigned( 215, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 831 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 30, 8)),
3 => std_logic_vector(to_unsigned( 142, 8)),
4 => std_logic_vector(to_unsigned( 133, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 45, 8)),
7 => std_logic_vector(to_unsigned( 235, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 159, 8)),
10 => std_logic_vector(to_unsigned( 32, 8)),
11 => std_logic_vector(to_unsigned( 248, 8)),
12 => std_logic_vector(to_unsigned( 147, 8)),
13 => std_logic_vector(to_unsigned( 134, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 153, 8)),
17 => std_logic_vector(to_unsigned( 178, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011101
elsif count = 832 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 212, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 212, 8)),
5 => std_logic_vector(to_unsigned( 87, 8)),
6 => std_logic_vector(to_unsigned( 122, 8)),
7 => std_logic_vector(to_unsigned( 247, 8)),
8 => std_logic_vector(to_unsigned( 209, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 128, 8)),
12 => std_logic_vector(to_unsigned( 153, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 90, 8)),
15 => std_logic_vector(to_unsigned( 185, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 159, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 833 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 161, 8)),
2 => std_logic_vector(to_unsigned( 101, 8)),
3 => std_logic_vector(to_unsigned( 59, 8)),
4 => std_logic_vector(to_unsigned( 65, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 123, 8)),
10 => std_logic_vector(to_unsigned( 1, 8)),
11 => std_logic_vector(to_unsigned( 120, 8)),
12 => std_logic_vector(to_unsigned( 136, 8)),
13 => std_logic_vector(to_unsigned( 190, 8)),
14 => std_logic_vector(to_unsigned( 68, 8)),
15 => std_logic_vector(to_unsigned( 72, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 123, 8)),
18 => std_logic_vector(to_unsigned( 70, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 834 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 142, 8)),
3 => std_logic_vector(to_unsigned( 50, 8)),
4 => std_logic_vector(to_unsigned( 75, 8)),
5 => std_logic_vector(to_unsigned( 88, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 246, 8)),
8 => std_logic_vector(to_unsigned( 31, 8)),
9 => std_logic_vector(to_unsigned( 70, 8)),
10 => std_logic_vector(to_unsigned( 127, 8)),
11 => std_logic_vector(to_unsigned( 107, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 232, 8)),
15 => std_logic_vector(to_unsigned( 130, 8)),
16 => std_logic_vector(to_unsigned( 49, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010101
elsif count = 835 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 169, 8)),
2 => std_logic_vector(to_unsigned( 162, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 141, 8)),
5 => std_logic_vector(to_unsigned( 9, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 94, 8)),
8 => std_logic_vector(to_unsigned( 240, 8)),
9 => std_logic_vector(to_unsigned( 237, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 59, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 43, 8)),
16 => std_logic_vector(to_unsigned( 215, 8)),
17 => std_logic_vector(to_unsigned( 52, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100110
elsif count = 836 then RAM <= (0 => "11111100",
1 => std_logic_vector(to_unsigned( 83, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 92, 8)),
5 => std_logic_vector(to_unsigned( 172, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 169, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 172, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 152, 8)),
12 => std_logic_vector(to_unsigned( 225, 8)),
13 => std_logic_vector(to_unsigned( 122, 8)),
14 => std_logic_vector(to_unsigned( 213, 8)),
15 => std_logic_vector(to_unsigned( 113, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 837 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 204, 8)),
2 => std_logic_vector(to_unsigned( 32, 8)),
3 => std_logic_vector(to_unsigned( 238, 8)),
4 => std_logic_vector(to_unsigned( 92, 8)),
5 => std_logic_vector(to_unsigned( 37, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 28, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 25, 8)),
11 => std_logic_vector(to_unsigned( 221, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 231, 8)),
15 => std_logic_vector(to_unsigned( 238, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110011
elsif count = 838 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 105, 8)),
2 => std_logic_vector(to_unsigned( 74, 8)),
3 => std_logic_vector(to_unsigned( 57, 8)),
4 => std_logic_vector(to_unsigned( 196, 8)),
5 => std_logic_vector(to_unsigned( 255, 8)),
6 => std_logic_vector(to_unsigned( 96, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 62, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 45, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 217, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 105, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 839 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 25, 8)),
2 => std_logic_vector(to_unsigned( 158, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 194, 8)),
5 => std_logic_vector(to_unsigned( 98, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 85, 8)),
8 => std_logic_vector(to_unsigned( 185, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 166, 8)),
11 => std_logic_vector(to_unsigned( 190, 8)),
12 => std_logic_vector(to_unsigned( 204, 8)),
13 => std_logic_vector(to_unsigned( 196, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 129, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 147, 8)),
18 => std_logic_vector(to_unsigned( 184, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 840 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 235, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 37, 8)),
5 => std_logic_vector(to_unsigned( 12, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 192, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 102, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 218, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 189, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 200, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 841 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 156, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 203, 8)),
4 => std_logic_vector(to_unsigned( 58, 8)),
5 => std_logic_vector(to_unsigned( 178, 8)),
6 => std_logic_vector(to_unsigned( 37, 8)),
7 => std_logic_vector(to_unsigned( 156, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 243, 8)),
10 => std_logic_vector(to_unsigned( 100, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 140, 8)),
13 => std_logic_vector(to_unsigned( 44, 8)),
14 => std_logic_vector(to_unsigned( 102, 8)),
15 => std_logic_vector(to_unsigned( 233, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 99, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 842 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 104, 8)),
3 => std_logic_vector(to_unsigned( 33, 8)),
4 => std_logic_vector(to_unsigned( 80, 8)),
5 => std_logic_vector(to_unsigned( 25, 8)),
6 => std_logic_vector(to_unsigned( 88, 8)),
7 => std_logic_vector(to_unsigned( 37, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 136, 8)),
11 => std_logic_vector(to_unsigned( 165, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 59, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 843 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 229, 8)),
2 => std_logic_vector(to_unsigned( 70, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 70, 8)),
8 => std_logic_vector(to_unsigned( 59, 8)),
9 => std_logic_vector(to_unsigned( 75, 8)),
10 => std_logic_vector(to_unsigned( 147, 8)),
11 => std_logic_vector(to_unsigned( 116, 8)),
12 => std_logic_vector(to_unsigned( 15, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 28, 8)),
15 => std_logic_vector(to_unsigned( 132, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 844 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 163, 8)),
4 => std_logic_vector(to_unsigned( 182, 8)),
5 => std_logic_vector(to_unsigned( 211, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 198, 8)),
8 => std_logic_vector(to_unsigned( 219, 8)),
9 => std_logic_vector(to_unsigned( 47, 8)),
10 => std_logic_vector(to_unsigned( 226, 8)),
11 => std_logic_vector(to_unsigned( 212, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 48, 8)),
14 => std_logic_vector(to_unsigned( 227, 8)),
15 => std_logic_vector(to_unsigned( 171, 8)),
16 => std_logic_vector(to_unsigned( 218, 8)),
17 => std_logic_vector(to_unsigned( 185, 8)),
18 => std_logic_vector(to_unsigned( 196, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101110
elsif count = 845 then RAM <= (0 => "01111110",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 44, 8)),
4 => std_logic_vector(to_unsigned( 77, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 119, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 68, 8)),
10 => std_logic_vector(to_unsigned( 121, 8)),
11 => std_logic_vector(to_unsigned( 46, 8)),
12 => std_logic_vector(to_unsigned( 101, 8)),
13 => std_logic_vector(to_unsigned( 68, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 6, 8)),
16 => std_logic_vector(to_unsigned( 97, 8)),
17 => std_logic_vector(to_unsigned( 67, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111110
elsif count = 846 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 131, 8)),
4 => std_logic_vector(to_unsigned( 55, 8)),
5 => std_logic_vector(to_unsigned( 68, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 98, 8)),
8 => std_logic_vector(to_unsigned( 159, 8)),
9 => std_logic_vector(to_unsigned( 77, 8)),
10 => std_logic_vector(to_unsigned( 33, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 177, 8)),
13 => std_logic_vector(to_unsigned( 183, 8)),
14 => std_logic_vector(to_unsigned( 199, 8)),
15 => std_logic_vector(to_unsigned( 131, 8)),
16 => std_logic_vector(to_unsigned( 29, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 42, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10010111
elsif count = 847 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 191, 8)),
2 => std_logic_vector(to_unsigned( 46, 8)),
3 => std_logic_vector(to_unsigned( 188, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 193, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 179, 8)),
8 => std_logic_vector(to_unsigned( 102, 8)),
9 => std_logic_vector(to_unsigned( 252, 8)),
10 => std_logic_vector(to_unsigned( 182, 8)),
11 => std_logic_vector(to_unsigned( 213, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 165, 8)),
14 => std_logic_vector(to_unsigned( 88, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 848 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 171, 8)),
2 => std_logic_vector(to_unsigned( 212, 8)),
3 => std_logic_vector(to_unsigned( 243, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 237, 8)),
7 => std_logic_vector(to_unsigned( 163, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 222, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 236, 8)),
13 => std_logic_vector(to_unsigned( 25, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 240, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 198, 8)),
18 => std_logic_vector(to_unsigned( 183, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 849 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 126, 8)),
3 => std_logic_vector(to_unsigned( 220, 8)),
4 => std_logic_vector(to_unsigned( 5, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 151, 8)),
7 => std_logic_vector(to_unsigned( 214, 8)),
8 => std_logic_vector(to_unsigned( 45, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 83, 8)),
11 => std_logic_vector(to_unsigned( 59, 8)),
12 => std_logic_vector(to_unsigned( 116, 8)),
13 => std_logic_vector(to_unsigned( 142, 8)),
14 => std_logic_vector(to_unsigned( 83, 8)),
15 => std_logic_vector(to_unsigned( 123, 8)),
16 => std_logic_vector(to_unsigned( 220, 8)),
17 => std_logic_vector(to_unsigned( 158, 8)),
18 => std_logic_vector(to_unsigned( 118, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 850 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 211, 8)),
2 => std_logic_vector(to_unsigned( 132, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 160, 8)),
5 => std_logic_vector(to_unsigned( 177, 8)),
6 => std_logic_vector(to_unsigned( 195, 8)),
7 => std_logic_vector(to_unsigned( 181, 8)),
8 => std_logic_vector(to_unsigned( 100, 8)),
9 => std_logic_vector(to_unsigned( 227, 8)),
10 => std_logic_vector(to_unsigned( 8, 8)),
11 => std_logic_vector(to_unsigned( 119, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 67, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 164, 8)),
16 => std_logic_vector(to_unsigned( 83, 8)),
17 => std_logic_vector(to_unsigned( 156, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 851 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 1, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 127, 8)),
4 => std_logic_vector(to_unsigned( 149, 8)),
5 => std_logic_vector(to_unsigned( 232, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 107, 8)),
9 => std_logic_vector(to_unsigned( 142, 8)),
10 => std_logic_vector(to_unsigned( 150, 8)),
11 => std_logic_vector(to_unsigned( 110, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 135, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 852 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 131, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 216, 8)),
4 => std_logic_vector(to_unsigned( 127, 8)),
5 => std_logic_vector(to_unsigned( 172, 8)),
6 => std_logic_vector(to_unsigned( 188, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 129, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 246, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 46, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 107, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 853 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 118, 8)),
3 => std_logic_vector(to_unsigned( 127, 8)),
4 => std_logic_vector(to_unsigned( 181, 8)),
5 => std_logic_vector(to_unsigned( 208, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 210, 8)),
8 => std_logic_vector(to_unsigned( 3, 8)),
9 => std_logic_vector(to_unsigned( 89, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 147, 8)),
12 => std_logic_vector(to_unsigned( 201, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 153, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 133, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 854 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 215, 8)),
2 => std_logic_vector(to_unsigned( 131, 8)),
3 => std_logic_vector(to_unsigned( 252, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 153, 8)),
6 => std_logic_vector(to_unsigned( 66, 8)),
7 => std_logic_vector(to_unsigned( 97, 8)),
8 => std_logic_vector(to_unsigned( 29, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 206, 8)),
12 => std_logic_vector(to_unsigned( 119, 8)),
13 => std_logic_vector(to_unsigned( 84, 8)),
14 => std_logic_vector(to_unsigned( 145, 8)),
15 => std_logic_vector(to_unsigned( 69, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 138, 8)),
18 => std_logic_vector(to_unsigned( 125, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110100
elsif count = 855 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 163, 8)),
2 => std_logic_vector(to_unsigned( 150, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 200, 8)),
6 => std_logic_vector(to_unsigned( 251, 8)),
7 => std_logic_vector(to_unsigned( 1, 8)),
8 => std_logic_vector(to_unsigned( 26, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 45, 8)),
11 => std_logic_vector(to_unsigned( 228, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 79, 8)),
14 => std_logic_vector(to_unsigned( 103, 8)),
15 => std_logic_vector(to_unsigned( 121, 8)),
16 => std_logic_vector(to_unsigned( 41, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 856 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 230, 8)),
2 => std_logic_vector(to_unsigned( 12, 8)),
3 => std_logic_vector(to_unsigned( 144, 8)),
4 => std_logic_vector(to_unsigned( 89, 8)),
5 => std_logic_vector(to_unsigned( 7, 8)),
6 => std_logic_vector(to_unsigned( 24, 8)),
7 => std_logic_vector(to_unsigned( 104, 8)),
8 => std_logic_vector(to_unsigned( 63, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 62, 8)),
11 => std_logic_vector(to_unsigned( 83, 8)),
12 => std_logic_vector(to_unsigned( 90, 8)),
13 => std_logic_vector(to_unsigned( 98, 8)),
14 => std_logic_vector(to_unsigned( 105, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 236, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 857 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 75, 8)),
2 => std_logic_vector(to_unsigned( 29, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 152, 8)),
5 => std_logic_vector(to_unsigned( 59, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 23, 8)),
9 => std_logic_vector(to_unsigned( 57, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 133, 8)),
13 => std_logic_vector(to_unsigned( 29, 8)),
14 => std_logic_vector(to_unsigned( 132, 8)),
15 => std_logic_vector(to_unsigned( 19, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 68, 8)),
18 => std_logic_vector(to_unsigned( 149, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 858 then RAM <= (0 => "11011110",
1 => std_logic_vector(to_unsigned( 70, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 255, 8)),
4 => std_logic_vector(to_unsigned( 142, 8)),
5 => std_logic_vector(to_unsigned( 22, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 65, 8)),
8 => std_logic_vector(to_unsigned( 78, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 18, 8)),
12 => std_logic_vector(to_unsigned( 156, 8)),
13 => std_logic_vector(to_unsigned( 87, 8)),
14 => std_logic_vector(to_unsigned( 112, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011000
elsif count = 859 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 134, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 140, 8)),
4 => std_logic_vector(to_unsigned( 8, 8)),
5 => std_logic_vector(to_unsigned( 214, 8)),
6 => std_logic_vector(to_unsigned( 203, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 172, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 75, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 26, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 89, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 86, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 69, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 860 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 84, 8)),
2 => std_logic_vector(to_unsigned( 34, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 34, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 233, 8)),
8 => std_logic_vector(to_unsigned( 230, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 207, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 86, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 95, 8)),
15 => std_logic_vector(to_unsigned( 63, 8)),
16 => std_logic_vector(to_unsigned( 43, 8)),
17 => std_logic_vector(to_unsigned( 110, 8)),
18 => std_logic_vector(to_unsigned( 55, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100110
elsif count = 861 then RAM <= (0 => "10111011",
1 => std_logic_vector(to_unsigned( 188, 8)),
2 => std_logic_vector(to_unsigned( 165, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 212, 8)),
5 => std_logic_vector(to_unsigned( 244, 8)),
6 => std_logic_vector(to_unsigned( 253, 8)),
7 => std_logic_vector(to_unsigned( 80, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 184, 8)),
11 => std_logic_vector(to_unsigned( 159, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 246, 8)),
15 => std_logic_vector(to_unsigned( 132, 8)),
16 => std_logic_vector(to_unsigned( 81, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111011
elsif count = 862 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 216, 8)),
5 => std_logic_vector(to_unsigned( 240, 8)),
6 => std_logic_vector(to_unsigned( 63, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 226, 8)),
9 => std_logic_vector(to_unsigned( 52, 8)),
10 => std_logic_vector(to_unsigned( 236, 8)),
11 => std_logic_vector(to_unsigned( 41, 8)),
12 => std_logic_vector(to_unsigned( 217, 8)),
13 => std_logic_vector(to_unsigned( 53, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 13, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 157, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 863 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 179, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 80, 8)),
5 => std_logic_vector(to_unsigned( 68, 8)),
6 => std_logic_vector(to_unsigned( 130, 8)),
7 => std_logic_vector(to_unsigned( 14, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 154, 8)),
11 => std_logic_vector(to_unsigned( 69, 8)),
12 => std_logic_vector(to_unsigned( 178, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 194, 8)),
15 => std_logic_vector(to_unsigned( 99, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 864 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 16, 8)),
4 => std_logic_vector(to_unsigned( 53, 8)),
5 => std_logic_vector(to_unsigned( 30, 8)),
6 => std_logic_vector(to_unsigned( 39, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 24, 8)),
10 => std_logic_vector(to_unsigned( 45, 8)),
11 => std_logic_vector(to_unsigned( 64, 8)),
12 => std_logic_vector(to_unsigned( 33, 8)),
13 => std_logic_vector(to_unsigned( 48, 8)),
14 => std_logic_vector(to_unsigned( 198, 8)),
15 => std_logic_vector(to_unsigned( 214, 8)),
16 => std_logic_vector(to_unsigned( 100, 8)),
17 => std_logic_vector(to_unsigned( 50, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110111
elsif count = 865 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 36, 8)),
3 => std_logic_vector(to_unsigned( 219, 8)),
4 => std_logic_vector(to_unsigned( 210, 8)),
5 => std_logic_vector(to_unsigned( 16, 8)),
6 => std_logic_vector(to_unsigned( 26, 8)),
7 => std_logic_vector(to_unsigned( 107, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 178, 8)),
10 => std_logic_vector(to_unsigned( 212, 8)),
11 => std_logic_vector(to_unsigned( 79, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 137, 8)),
16 => std_logic_vector(to_unsigned( 32, 8)),
17 => std_logic_vector(to_unsigned( 124, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 866 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 192, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 61, 8)),
5 => std_logic_vector(to_unsigned( 53, 8)),
6 => std_logic_vector(to_unsigned( 235, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 18, 8)),
10 => std_logic_vector(to_unsigned( 214, 8)),
11 => std_logic_vector(to_unsigned( 23, 8)),
12 => std_logic_vector(to_unsigned( 113, 8)),
13 => std_logic_vector(to_unsigned( 22, 8)),
14 => std_logic_vector(to_unsigned( 114, 8)),
15 => std_logic_vector(to_unsigned( 195, 8)),
16 => std_logic_vector(to_unsigned( 177, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 867 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 244, 8)),
2 => std_logic_vector(to_unsigned( 41, 8)),
3 => std_logic_vector(to_unsigned( 55, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 97, 8)),
6 => std_logic_vector(to_unsigned( 179, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 223, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 157, 8)),
12 => std_logic_vector(to_unsigned( 210, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 160, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 868 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 44, 8)),
3 => std_logic_vector(to_unsigned( 62, 8)),
4 => std_logic_vector(to_unsigned( 15, 8)),
5 => std_logic_vector(to_unsigned( 76, 8)),
6 => std_logic_vector(to_unsigned( 149, 8)),
7 => std_logic_vector(to_unsigned( 49, 8)),
8 => std_logic_vector(to_unsigned( 28, 8)),
9 => std_logic_vector(to_unsigned( 120, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 164, 8)),
12 => std_logic_vector(to_unsigned( 237, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 213, 8)),
15 => std_logic_vector(to_unsigned( 33, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 869 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 66, 8)),
2 => std_logic_vector(to_unsigned( 136, 8)),
3 => std_logic_vector(to_unsigned( 108, 8)),
4 => std_logic_vector(to_unsigned( 94, 8)),
5 => std_logic_vector(to_unsigned( 208, 8)),
6 => std_logic_vector(to_unsigned( 115, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 190, 8)),
9 => std_logic_vector(to_unsigned( 13, 8)),
10 => std_logic_vector(to_unsigned( 243, 8)),
11 => std_logic_vector(to_unsigned( 93, 8)),
12 => std_logic_vector(to_unsigned( 109, 8)),
13 => std_logic_vector(to_unsigned( 140, 8)),
14 => std_logic_vector(to_unsigned( 172, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 190, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 870 then RAM <= (0 => "11110011",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 64, 8)),
3 => std_logic_vector(to_unsigned( 168, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 29, 8)),
7 => std_logic_vector(to_unsigned( 193, 8)),
8 => std_logic_vector(to_unsigned( 19, 8)),
9 => std_logic_vector(to_unsigned( 83, 8)),
10 => std_logic_vector(to_unsigned( 175, 8)),
11 => std_logic_vector(to_unsigned( 114, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 118, 8)),
14 => std_logic_vector(to_unsigned( 216, 8)),
15 => std_logic_vector(to_unsigned( 50, 8)),
16 => std_logic_vector(to_unsigned( 250, 8)),
17 => std_logic_vector(to_unsigned( 152, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 871 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 166, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 116, 8)),
6 => std_logic_vector(to_unsigned( 79, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 112, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 155, 8)),
13 => std_logic_vector(to_unsigned( 249, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 144, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 126, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 872 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 142, 8)),
2 => std_logic_vector(to_unsigned( 249, 8)),
3 => std_logic_vector(to_unsigned( 127, 8)),
4 => std_logic_vector(to_unsigned( 77, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 152, 8)),
7 => std_logic_vector(to_unsigned( 211, 8)),
8 => std_logic_vector(to_unsigned( 135, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 245, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 252, 8)),
13 => std_logic_vector(to_unsigned( 100, 8)),
14 => std_logic_vector(to_unsigned( 104, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 177, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 143, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001110
elsif count = 873 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 147, 8)),
2 => std_logic_vector(to_unsigned( 202, 8)),
3 => std_logic_vector(to_unsigned( 146, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 18, 8)),
6 => std_logic_vector(to_unsigned( 175, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 105, 8)),
9 => std_logic_vector(to_unsigned( 254, 8)),
10 => std_logic_vector(to_unsigned( 7, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 223, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 114, 8)),
16 => std_logic_vector(to_unsigned( 27, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01100111
elsif count = 874 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 44, 8)),
5 => std_logic_vector(to_unsigned( 201, 8)),
6 => std_logic_vector(to_unsigned( 58, 8)),
7 => std_logic_vector(to_unsigned( 30, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 57, 8)),
11 => std_logic_vector(to_unsigned( 242, 8)),
12 => std_logic_vector(to_unsigned( 10, 8)),
13 => std_logic_vector(to_unsigned( 211, 8)),
14 => std_logic_vector(to_unsigned( 76, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 58, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 72, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 875 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 33, 8)),
3 => std_logic_vector(to_unsigned( 178, 8)),
4 => std_logic_vector(to_unsigned( 112, 8)),
5 => std_logic_vector(to_unsigned( 206, 8)),
6 => std_logic_vector(to_unsigned( 32, 8)),
7 => std_logic_vector(to_unsigned( 181, 8)),
8 => std_logic_vector(to_unsigned( 39, 8)),
9 => std_logic_vector(to_unsigned( 44, 8)),
10 => std_logic_vector(to_unsigned( 213, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 81, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 102, 8)),
17 => std_logic_vector(to_unsigned( 144, 8)),
18 => std_logic_vector(to_unsigned( 65, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101001
elsif count = 876 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 189, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 208, 8)),
5 => std_logic_vector(to_unsigned( 156, 8)),
6 => std_logic_vector(to_unsigned( 51, 8)),
7 => std_logic_vector(to_unsigned( 223, 8)),
8 => std_logic_vector(to_unsigned( 148, 8)),
9 => std_logic_vector(to_unsigned( 115, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 103, 8)),
12 => std_logic_vector(to_unsigned( 205, 8)),
13 => std_logic_vector(to_unsigned( 42, 8)),
14 => std_logic_vector(to_unsigned( 190, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 41, 8)),
17 => std_logic_vector(to_unsigned( 80, 8)),
18 => std_logic_vector(to_unsigned( 187, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 877 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 58, 8)),
3 => std_logic_vector(to_unsigned( 70, 8)),
4 => std_logic_vector(to_unsigned( 140, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 206, 8)),
7 => std_logic_vector(to_unsigned( 91, 8)),
8 => std_logic_vector(to_unsigned( 71, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 51, 8)),
11 => std_logic_vector(to_unsigned( 203, 8)),
12 => std_logic_vector(to_unsigned( 248, 8)),
13 => std_logic_vector(to_unsigned( 129, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 62, 8)),
17 => std_logic_vector(to_unsigned( 121, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 878 then RAM <= (0 => "01110111",
1 => std_logic_vector(to_unsigned( 152, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 151, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 163, 8)),
6 => std_logic_vector(to_unsigned( 111, 8)),
7 => std_logic_vector(to_unsigned( 227, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 85, 8)),
10 => std_logic_vector(to_unsigned( 244, 8)),
11 => std_logic_vector(to_unsigned( 170, 8)),
12 => std_logic_vector(to_unsigned( 61, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 49, 8)),
15 => std_logic_vector(to_unsigned( 254, 8)),
16 => std_logic_vector(to_unsigned( 36, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01000111
elsif count = 879 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 112, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 63, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 95, 8)),
10 => std_logic_vector(to_unsigned( 205, 8)),
11 => std_logic_vector(to_unsigned( 36, 8)),
12 => std_logic_vector(to_unsigned( 220, 8)),
13 => std_logic_vector(to_unsigned( 113, 8)),
14 => std_logic_vector(to_unsigned( 187, 8)),
15 => std_logic_vector(to_unsigned( 219, 8)),
16 => std_logic_vector(to_unsigned( 255, 8)),
17 => std_logic_vector(to_unsigned( 58, 8)),
18 => std_logic_vector(to_unsigned( 187, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111001
elsif count = 880 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 187, 8)),
2 => std_logic_vector(to_unsigned( 151, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 54, 8)),
5 => std_logic_vector(to_unsigned( 172, 8)),
6 => std_logic_vector(to_unsigned( 106, 8)),
7 => std_logic_vector(to_unsigned( 88, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 84, 8)),
11 => std_logic_vector(to_unsigned( 180, 8)),
12 => std_logic_vector(to_unsigned( 114, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 110, 8)),
15 => std_logic_vector(to_unsigned( 83, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 119, 8)),
18 => std_logic_vector(to_unsigned( 126, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 881 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 200, 8)),
3 => std_logic_vector(to_unsigned( 156, 8)),
4 => std_logic_vector(to_unsigned( 75, 8)),
5 => std_logic_vector(to_unsigned( 175, 8)),
6 => std_logic_vector(to_unsigned( 231, 8)),
7 => std_logic_vector(to_unsigned( 187, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 30, 8)),
10 => std_logic_vector(to_unsigned( 77, 8)),
11 => std_logic_vector(to_unsigned( 191, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 199, 8)),
14 => std_logic_vector(to_unsigned( 229, 8)),
15 => std_logic_vector(to_unsigned( 170, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 186, 8)),
18 => std_logic_vector(to_unsigned( 193, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 882 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 145, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 19, 8)),
5 => std_logic_vector(to_unsigned( 224, 8)),
6 => std_logic_vector(to_unsigned( 55, 8)),
7 => std_logic_vector(to_unsigned( 76, 8)),
8 => std_logic_vector(to_unsigned( 177, 8)),
9 => std_logic_vector(to_unsigned( 147, 8)),
10 => std_logic_vector(to_unsigned( 120, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 136, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 98, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 116, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111000
elsif count = 883 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 36, 8)),
2 => std_logic_vector(to_unsigned( 118, 8)),
3 => std_logic_vector(to_unsigned( 211, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 157, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 125, 8)),
9 => std_logic_vector(to_unsigned( 171, 8)),
10 => std_logic_vector(to_unsigned( 133, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 130, 8)),
13 => std_logic_vector(to_unsigned( 144, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 163, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110110
elsif count = 884 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 213, 8)),
2 => std_logic_vector(to_unsigned( 135, 8)),
3 => std_logic_vector(to_unsigned( 200, 8)),
4 => std_logic_vector(to_unsigned( 140, 8)),
5 => std_logic_vector(to_unsigned( 35, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 149, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 167, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 87, 8)),
15 => std_logic_vector(to_unsigned( 140, 8)),
16 => std_logic_vector(to_unsigned( 200, 8)),
17 => std_logic_vector(to_unsigned( 131, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 885 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 140, 8)),
3 => std_logic_vector(to_unsigned( 45, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 24, 8)),
6 => std_logic_vector(to_unsigned( 178, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 49, 8)),
10 => std_logic_vector(to_unsigned( 186, 8)),
11 => std_logic_vector(to_unsigned( 55, 8)),
12 => std_logic_vector(to_unsigned( 199, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 100, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 134, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 886 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 70, 8)),
5 => std_logic_vector(to_unsigned( 35, 8)),
6 => std_logic_vector(to_unsigned( 7, 8)),
7 => std_logic_vector(to_unsigned( 66, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 113, 8)),
10 => std_logic_vector(to_unsigned( 79, 8)),
11 => std_logic_vector(to_unsigned( 39, 8)),
12 => std_logic_vector(to_unsigned( 247, 8)),
13 => std_logic_vector(to_unsigned( 155, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 149, 8)),
16 => std_logic_vector(to_unsigned( 133, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 124, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 887 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 184, 8)),
2 => std_logic_vector(to_unsigned( 169, 8)),
3 => std_logic_vector(to_unsigned( 213, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 165, 8)),
7 => std_logic_vector(to_unsigned( 87, 8)),
8 => std_logic_vector(to_unsigned( 174, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 98, 8)),
11 => std_logic_vector(to_unsigned( 181, 8)),
12 => std_logic_vector(to_unsigned( 172, 8)),
13 => std_logic_vector(to_unsigned( 234, 8)),
14 => std_logic_vector(to_unsigned( 183, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 192, 8)),
17 => std_logic_vector(to_unsigned( 202, 8)),
18 => std_logic_vector(to_unsigned( 195, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 888 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 135, 8)),
2 => std_logic_vector(to_unsigned( 209, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 247, 8)),
5 => std_logic_vector(to_unsigned( 182, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 153, 8)),
8 => std_logic_vector(to_unsigned( 66, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 69, 8)),
11 => std_logic_vector(to_unsigned( 210, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 254, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111100
elsif count = 889 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 77, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 167, 8)),
5 => std_logic_vector(to_unsigned( 83, 8)),
6 => std_logic_vector(to_unsigned( 170, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 133, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 229, 8)),
12 => std_logic_vector(to_unsigned( 60, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 162, 8)),
16 => std_logic_vector(to_unsigned( 74, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 134, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 890 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 11, 8)),
2 => std_logic_vector(to_unsigned( 205, 8)),
3 => std_logic_vector(to_unsigned( 164, 8)),
4 => std_logic_vector(to_unsigned( 219, 8)),
5 => std_logic_vector(to_unsigned( 3, 8)),
6 => std_logic_vector(to_unsigned( 230, 8)),
7 => std_logic_vector(to_unsigned( 190, 8)),
8 => std_logic_vector(to_unsigned( 245, 8)),
9 => std_logic_vector(to_unsigned( 204, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 148, 8)),
12 => std_logic_vector(to_unsigned( 181, 8)),
13 => std_logic_vector(to_unsigned( 217, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 54, 8)),
16 => std_logic_vector(to_unsigned( 176, 8)),
17 => std_logic_vector(to_unsigned( 191, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111010
elsif count = 891 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 223, 8)),
2 => std_logic_vector(to_unsigned( 99, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 162, 8)),
5 => std_logic_vector(to_unsigned( 79, 8)),
6 => std_logic_vector(to_unsigned( 56, 8)),
7 => std_logic_vector(to_unsigned( 144, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 197, 8)),
10 => std_logic_vector(to_unsigned( 193, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 69, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 44, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 121, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001100
elsif count = 892 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 0, 8)),
4 => std_logic_vector(to_unsigned( 89, 8)),
5 => std_logic_vector(to_unsigned( 20, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 48, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 82, 8)),
10 => std_logic_vector(to_unsigned( 24, 8)),
11 => std_logic_vector(to_unsigned( 88, 8)),
12 => std_logic_vector(to_unsigned( 55, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 63, 8)),
15 => std_logic_vector(to_unsigned( 34, 8)),
16 => std_logic_vector(to_unsigned( 99, 8)),
17 => std_logic_vector(to_unsigned( 64, 8)),
18 => std_logic_vector(to_unsigned( 80, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 893 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 233, 8)),
4 => std_logic_vector(to_unsigned( 176, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 142, 8)),
7 => std_logic_vector(to_unsigned( 186, 8)),
8 => std_logic_vector(to_unsigned( 11, 8)),
9 => std_logic_vector(to_unsigned( 48, 8)),
10 => std_logic_vector(to_unsigned( 66, 8)),
11 => std_logic_vector(to_unsigned( 215, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 106, 8)),
14 => std_logic_vector(to_unsigned( 72, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 74, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 894 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 245, 8)),
2 => std_logic_vector(to_unsigned( 89, 8)),
3 => std_logic_vector(to_unsigned( 58, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 48, 8)),
7 => std_logic_vector(to_unsigned( 146, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 79, 8)),
10 => std_logic_vector(to_unsigned( 21, 8)),
11 => std_logic_vector(to_unsigned( 91, 8)),
12 => std_logic_vector(to_unsigned( 11, 8)),
13 => std_logic_vector(to_unsigned( 63, 8)),
14 => std_logic_vector(to_unsigned( 39, 8)),
15 => std_logic_vector(to_unsigned( 14, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 100, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101100
elsif count = 895 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 143, 8)),
2 => std_logic_vector(to_unsigned( 116, 8)),
3 => std_logic_vector(to_unsigned( 91, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 130, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 13, 8)),
8 => std_logic_vector(to_unsigned( 55, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 12, 8)),
11 => std_logic_vector(to_unsigned( 108, 8)),
12 => std_logic_vector(to_unsigned( 171, 8)),
13 => std_logic_vector(to_unsigned( 56, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 97, 8)),
16 => std_logic_vector(to_unsigned( 98, 8)),
17 => std_logic_vector(to_unsigned( 111, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 896 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 110, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 175, 8)),
4 => std_logic_vector(to_unsigned( 161, 8)),
5 => std_logic_vector(to_unsigned( 217, 8)),
6 => std_logic_vector(to_unsigned( 92, 8)),
7 => std_logic_vector(to_unsigned( 59, 8)),
8 => std_logic_vector(to_unsigned( 88, 8)),
9 => std_logic_vector(to_unsigned( 135, 8)),
10 => std_logic_vector(to_unsigned( 97, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 114, 8)),
14 => std_logic_vector(to_unsigned( 118, 8)),
15 => std_logic_vector(to_unsigned( 156, 8)),
16 => std_logic_vector(to_unsigned( 180, 8)),
17 => std_logic_vector(to_unsigned( 140, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 897 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 49, 8)),
3 => std_logic_vector(to_unsigned( 37, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 65, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 57, 8)),
8 => std_logic_vector(to_unsigned( 147, 8)),
9 => std_logic_vector(to_unsigned( 128, 8)),
10 => std_logic_vector(to_unsigned( 94, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 115, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 151, 8)),
15 => std_logic_vector(to_unsigned( 62, 8)),
16 => std_logic_vector(to_unsigned( 70, 8)),
17 => std_logic_vector(to_unsigned( 61, 8)),
18 => std_logic_vector(to_unsigned( 110, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101110
elsif count = 898 then RAM <= (0 => "01011111",
1 => std_logic_vector(to_unsigned( 216, 8)),
2 => std_logic_vector(to_unsigned( 186, 8)),
3 => std_logic_vector(to_unsigned( 228, 8)),
4 => std_logic_vector(to_unsigned( 172, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 192, 8)),
7 => std_logic_vector(to_unsigned( 201, 8)),
8 => std_logic_vector(to_unsigned( 145, 8)),
9 => std_logic_vector(to_unsigned( 151, 8)),
10 => std_logic_vector(to_unsigned( 129, 8)),
11 => std_logic_vector(to_unsigned( 215, 8)),
12 => std_logic_vector(to_unsigned( 236, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 209, 8)),
15 => std_logic_vector(to_unsigned( 113, 8)),
16 => std_logic_vector(to_unsigned( 189, 8)),
17 => std_logic_vector(to_unsigned( 168, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011111
elsif count = 899 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 62, 8)),
3 => std_logic_vector(to_unsigned( 126, 8)),
4 => std_logic_vector(to_unsigned( 5, 8)),
5 => std_logic_vector(to_unsigned( 196, 8)),
6 => std_logic_vector(to_unsigned( 100, 8)),
7 => std_logic_vector(to_unsigned( 12, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 115, 8)),
11 => std_logic_vector(to_unsigned( 218, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 203, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 182, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000101
elsif count = 900 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 79, 8)),
3 => std_logic_vector(to_unsigned( 233, 8)),
4 => std_logic_vector(to_unsigned( 241, 8)),
5 => std_logic_vector(to_unsigned( 30, 8)),
6 => std_logic_vector(to_unsigned( 91, 8)),
7 => std_logic_vector(to_unsigned( 226, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 48, 8)),
10 => std_logic_vector(to_unsigned( 43, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 48, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 65, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 59, 8)),
18 => std_logic_vector(to_unsigned( 76, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010101
elsif count = 901 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 53, 8)),
2 => std_logic_vector(to_unsigned( 123, 8)),
3 => std_logic_vector(to_unsigned( 72, 8)),
4 => std_logic_vector(to_unsigned( 104, 8)),
5 => std_logic_vector(to_unsigned( 168, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 52, 8)),
8 => std_logic_vector(to_unsigned( 188, 8)),
9 => std_logic_vector(to_unsigned( 186, 8)),
10 => std_logic_vector(to_unsigned( 88, 8)),
11 => std_logic_vector(to_unsigned( 100, 8)),
12 => std_logic_vector(to_unsigned( 96, 8)),
13 => std_logic_vector(to_unsigned( 22, 8)),
14 => std_logic_vector(to_unsigned( 51, 8)),
15 => std_logic_vector(to_unsigned( 141, 8)),
16 => std_logic_vector(to_unsigned( 137, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100011
elsif count = 902 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 215, 8)),
2 => std_logic_vector(to_unsigned( 148, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 144, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 147, 8)),
7 => std_logic_vector(to_unsigned( 151, 8)),
8 => std_logic_vector(to_unsigned( 240, 8)),
9 => std_logic_vector(to_unsigned( 45, 8)),
10 => std_logic_vector(to_unsigned( 99, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 228, 8)),
13 => std_logic_vector(to_unsigned( 196, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 236, 8)),
16 => std_logic_vector(to_unsigned( 169, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100111
elsif count = 903 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 170, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 48, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 40, 8)),
7 => std_logic_vector(to_unsigned( 58, 8)),
8 => std_logic_vector(to_unsigned( 130, 8)),
9 => std_logic_vector(to_unsigned( 164, 8)),
10 => std_logic_vector(to_unsigned( 37, 8)),
11 => std_logic_vector(to_unsigned( 166, 8)),
12 => std_logic_vector(to_unsigned( 79, 8)),
13 => std_logic_vector(to_unsigned( 164, 8)),
14 => std_logic_vector(to_unsigned( 81, 8)),
15 => std_logic_vector(to_unsigned( 132, 8)),
16 => std_logic_vector(to_unsigned( 33, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 904 then RAM <= (0 => "10111101",
1 => std_logic_vector(to_unsigned( 236, 8)),
2 => std_logic_vector(to_unsigned( 163, 8)),
3 => std_logic_vector(to_unsigned( 201, 8)),
4 => std_logic_vector(to_unsigned( 236, 8)),
5 => std_logic_vector(to_unsigned( 221, 8)),
6 => std_logic_vector(to_unsigned( 200, 8)),
7 => std_logic_vector(to_unsigned( 226, 8)),
8 => std_logic_vector(to_unsigned( 153, 8)),
9 => std_logic_vector(to_unsigned( 116, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 237, 8)),
12 => std_logic_vector(to_unsigned( 184, 8)),
13 => std_logic_vector(to_unsigned( 128, 8)),
14 => std_logic_vector(to_unsigned( 215, 8)),
15 => std_logic_vector(to_unsigned( 106, 8)),
16 => std_logic_vector(to_unsigned( 178, 8)),
17 => std_logic_vector(to_unsigned( 203, 8)),
18 => std_logic_vector(to_unsigned( 174, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 905 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 166, 8)),
3 => std_logic_vector(to_unsigned( 183, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 239, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 57, 8)),
8 => std_logic_vector(to_unsigned( 67, 8)),
9 => std_logic_vector(to_unsigned( 17, 8)),
10 => std_logic_vector(to_unsigned( 91, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 227, 8)),
13 => std_logic_vector(to_unsigned( 210, 8)),
14 => std_logic_vector(to_unsigned( 93, 8)),
15 => std_logic_vector(to_unsigned( 224, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 193, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000111
elsif count = 906 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 98, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 126, 8)),
6 => std_logic_vector(to_unsigned( 109, 8)),
7 => std_logic_vector(to_unsigned( 249, 8)),
8 => std_logic_vector(to_unsigned( 164, 8)),
9 => std_logic_vector(to_unsigned( 105, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 138, 8)),
12 => std_logic_vector(to_unsigned( 57, 8)),
13 => std_logic_vector(to_unsigned( 30, 8)),
14 => std_logic_vector(to_unsigned( 166, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 93, 8)),
17 => std_logic_vector(to_unsigned( 115, 8)),
18 => std_logic_vector(to_unsigned( 77, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 907 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 107, 8)),
2 => std_logic_vector(to_unsigned( 19, 8)),
3 => std_logic_vector(to_unsigned( 114, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 75, 8)),
6 => std_logic_vector(to_unsigned( 190, 8)),
7 => std_logic_vector(to_unsigned( 114, 8)),
8 => std_logic_vector(to_unsigned( 237, 8)),
9 => std_logic_vector(to_unsigned( 73, 8)),
10 => std_logic_vector(to_unsigned( 192, 8)),
11 => std_logic_vector(to_unsigned( 95, 8)),
12 => std_logic_vector(to_unsigned( 170, 8)),
13 => std_logic_vector(to_unsigned( 76, 8)),
14 => std_logic_vector(to_unsigned( 177, 8)),
15 => std_logic_vector(to_unsigned( 173, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 194, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 908 then RAM <= (0 => "11011101",
1 => std_logic_vector(to_unsigned( 124, 8)),
2 => std_logic_vector(to_unsigned( 180, 8)),
3 => std_logic_vector(to_unsigned( 206, 8)),
4 => std_logic_vector(to_unsigned( 224, 8)),
5 => std_logic_vector(to_unsigned( 47, 8)),
6 => std_logic_vector(to_unsigned( 176, 8)),
7 => std_logic_vector(to_unsigned( 92, 8)),
8 => std_logic_vector(to_unsigned( 110, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 190, 8)),
11 => std_logic_vector(to_unsigned( 227, 8)),
12 => std_logic_vector(to_unsigned( 139, 8)),
13 => std_logic_vector(to_unsigned( 82, 8)),
14 => std_logic_vector(to_unsigned( 138, 8)),
15 => std_logic_vector(to_unsigned( 20, 8)),
16 => std_logic_vector(to_unsigned( 107, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 129, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011001
elsif count = 909 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 183, 8)),
2 => std_logic_vector(to_unsigned( 50, 8)),
3 => std_logic_vector(to_unsigned( 170, 8)),
4 => std_logic_vector(to_unsigned( 143, 8)),
5 => std_logic_vector(to_unsigned( 226, 8)),
6 => std_logic_vector(to_unsigned( 93, 8)),
7 => std_logic_vector(to_unsigned( 210, 8)),
8 => std_logic_vector(to_unsigned( 141, 8)),
9 => std_logic_vector(to_unsigned( 65, 8)),
10 => std_logic_vector(to_unsigned( 251, 8)),
11 => std_logic_vector(to_unsigned( 173, 8)),
12 => std_logic_vector(to_unsigned( 146, 8)),
13 => std_logic_vector(to_unsigned( 251, 8)),
14 => std_logic_vector(to_unsigned( 117, 8)),
15 => std_logic_vector(to_unsigned( 222, 8)),
16 => std_logic_vector(to_unsigned( 162, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 95, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00100111
elsif count = 910 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 205, 8)),
2 => std_logic_vector(to_unsigned( 199, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 131, 8)),
5 => std_logic_vector(to_unsigned( 122, 8)),
6 => std_logic_vector(to_unsigned( 177, 8)),
7 => std_logic_vector(to_unsigned( 69, 8)),
8 => std_logic_vector(to_unsigned( 230, 8)),
9 => std_logic_vector(to_unsigned( 22, 8)),
10 => std_logic_vector(to_unsigned( 159, 8)),
11 => std_logic_vector(to_unsigned( 141, 8)),
12 => std_logic_vector(to_unsigned( 194, 8)),
13 => std_logic_vector(to_unsigned( 39, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 41, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 69, 8)),
18 => std_logic_vector(to_unsigned( 171, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011110
elsif count = 911 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 116, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 98, 8)),
4 => std_logic_vector(to_unsigned( 137, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 203, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 204, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 41, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 213, 8)),
14 => std_logic_vector(to_unsigned( 65, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 91, 8)),
18 => std_logic_vector(to_unsigned( 88, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10000111
elsif count = 912 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 63, 8)),
2 => std_logic_vector(to_unsigned( 139, 8)),
3 => std_logic_vector(to_unsigned( 140, 8)),
4 => std_logic_vector(to_unsigned( 84, 8)),
5 => std_logic_vector(to_unsigned( 180, 8)),
6 => std_logic_vector(to_unsigned( 103, 8)),
7 => std_logic_vector(to_unsigned( 122, 8)),
8 => std_logic_vector(to_unsigned( 66, 8)),
9 => std_logic_vector(to_unsigned( 60, 8)),
10 => std_logic_vector(to_unsigned( 35, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 66, 8)),
13 => std_logic_vector(to_unsigned( 112, 8)),
14 => std_logic_vector(to_unsigned( 196, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 151, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 87, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101011
elsif count = 913 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 201, 8)),
2 => std_logic_vector(to_unsigned( 196, 8)),
3 => std_logic_vector(to_unsigned( 161, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 172, 8)),
7 => std_logic_vector(to_unsigned( 155, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 131, 8)),
10 => std_logic_vector(to_unsigned( 184, 8)),
11 => std_logic_vector(to_unsigned( 95, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 59, 8)),
14 => std_logic_vector(to_unsigned( 142, 8)),
15 => std_logic_vector(to_unsigned( 78, 8)),
16 => std_logic_vector(to_unsigned( 123, 8)),
17 => std_logic_vector(to_unsigned( 116, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 914 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 240, 8)),
2 => std_logic_vector(to_unsigned( 229, 8)),
3 => std_logic_vector(to_unsigned( 213, 8)),
4 => std_logic_vector(to_unsigned( 189, 8)),
5 => std_logic_vector(to_unsigned( 151, 8)),
6 => std_logic_vector(to_unsigned( 197, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 128, 8)),
9 => std_logic_vector(to_unsigned( 106, 8)),
10 => std_logic_vector(to_unsigned( 190, 8)),
11 => std_logic_vector(to_unsigned( 73, 8)),
12 => std_logic_vector(to_unsigned( 179, 8)),
13 => std_logic_vector(to_unsigned( 224, 8)),
14 => std_logic_vector(to_unsigned( 48, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 194, 8)),
17 => std_logic_vector(to_unsigned( 132, 8)),
18 => std_logic_vector(to_unsigned( 169, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011100
elsif count = 915 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 223, 8)),
2 => std_logic_vector(to_unsigned( 147, 8)),
3 => std_logic_vector(to_unsigned( 73, 8)),
4 => std_logic_vector(to_unsigned( 68, 8)),
5 => std_logic_vector(to_unsigned( 58, 8)),
6 => std_logic_vector(to_unsigned( 112, 8)),
7 => std_logic_vector(to_unsigned( 164, 8)),
8 => std_logic_vector(to_unsigned( 49, 8)),
9 => std_logic_vector(to_unsigned( 165, 8)),
10 => std_logic_vector(to_unsigned( 96, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 84, 8)),
13 => std_logic_vector(to_unsigned( 195, 8)),
14 => std_logic_vector(to_unsigned( 234, 8)),
15 => std_logic_vector(to_unsigned( 152, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 73, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111010
elsif count = 916 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 172, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 87, 8)),
4 => std_logic_vector(to_unsigned( 157, 8)),
5 => std_logic_vector(to_unsigned( 53, 8)),
6 => std_logic_vector(to_unsigned( 117, 8)),
7 => std_logic_vector(to_unsigned( 84, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 107, 8)),
10 => std_logic_vector(to_unsigned( 231, 8)),
11 => std_logic_vector(to_unsigned( 211, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 162, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 120, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 917 then RAM <= (0 => "11110101",
1 => std_logic_vector(to_unsigned( 43, 8)),
2 => std_logic_vector(to_unsigned( 149, 8)),
3 => std_logic_vector(to_unsigned( 253, 8)),
4 => std_logic_vector(to_unsigned( 111, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 67, 8)),
7 => std_logic_vector(to_unsigned( 165, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 109, 8)),
13 => std_logic_vector(to_unsigned( 94, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 109, 8)),
16 => std_logic_vector(to_unsigned( 63, 8)),
17 => std_logic_vector(to_unsigned( 105, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110101
elsif count = 918 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 70, 8)),
2 => std_logic_vector(to_unsigned( 230, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 80, 8)),
6 => std_logic_vector(to_unsigned( 220, 8)),
7 => std_logic_vector(to_unsigned( 7, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 117, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 201, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 215, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 42, 8)),
17 => std_logic_vector(to_unsigned( 62, 8)),
18 => std_logic_vector(to_unsigned( 182, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 919 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 199, 8)),
2 => std_logic_vector(to_unsigned( 67, 8)),
3 => std_logic_vector(to_unsigned( 205, 8)),
4 => std_logic_vector(to_unsigned( 69, 8)),
5 => std_logic_vector(to_unsigned( 40, 8)),
6 => std_logic_vector(to_unsigned( 196, 8)),
7 => std_logic_vector(to_unsigned( 244, 8)),
8 => std_logic_vector(to_unsigned( 98, 8)),
9 => std_logic_vector(to_unsigned( 42, 8)),
10 => std_logic_vector(to_unsigned( 37, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 215, 8)),
14 => std_logic_vector(to_unsigned( 79, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 92, 8)),
17 => std_logic_vector(to_unsigned( 201, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100011
elsif count = 920 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 181, 8)),
2 => std_logic_vector(to_unsigned( 86, 8)),
3 => std_logic_vector(to_unsigned( 194, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 40, 8)),
10 => std_logic_vector(to_unsigned( 31, 8)),
11 => std_logic_vector(to_unsigned( 99, 8)),
12 => std_logic_vector(to_unsigned( 221, 8)),
13 => std_logic_vector(to_unsigned( 87, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 94, 8)),
16 => std_logic_vector(to_unsigned( 130, 8)),
17 => std_logic_vector(to_unsigned( 90, 8)),
18 => std_logic_vector(to_unsigned( 178, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 921 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 122, 8)),
4 => std_logic_vector(to_unsigned( 222, 8)),
5 => std_logic_vector(to_unsigned( 233, 8)),
6 => std_logic_vector(to_unsigned( 34, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 41, 8)),
9 => std_logic_vector(to_unsigned( 220, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 154, 8)),
12 => std_logic_vector(to_unsigned( 231, 8)),
13 => std_logic_vector(to_unsigned( 116, 8)),
14 => std_logic_vector(to_unsigned( 159, 8)),
15 => std_logic_vector(to_unsigned( 159, 8)),
16 => std_logic_vector(to_unsigned( 116, 8)),
17 => std_logic_vector(to_unsigned( 176, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110000
elsif count = 922 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 30, 8)),
3 => std_logic_vector(to_unsigned( 212, 8)),
4 => std_logic_vector(to_unsigned( 139, 8)),
5 => std_logic_vector(to_unsigned( 150, 8)),
6 => std_logic_vector(to_unsigned( 198, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 187, 8)),
10 => std_logic_vector(to_unsigned( 195, 8)),
11 => std_logic_vector(to_unsigned( 189, 8)),
12 => std_logic_vector(to_unsigned( 223, 8)),
13 => std_logic_vector(to_unsigned( 148, 8)),
14 => std_logic_vector(to_unsigned( 200, 8)),
15 => std_logic_vector(to_unsigned( 180, 8)),
16 => std_logic_vector(to_unsigned( 232, 8)),
17 => std_logic_vector(to_unsigned( 170, 8)),
18 => std_logic_vector(to_unsigned( 210, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111100
elsif count = 923 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 185, 8)),
2 => std_logic_vector(to_unsigned( 24, 8)),
3 => std_logic_vector(to_unsigned( 77, 8)),
4 => std_logic_vector(to_unsigned( 87, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 22, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 195, 8)),
10 => std_logic_vector(to_unsigned( 134, 8)),
11 => std_logic_vector(to_unsigned( 42, 8)),
12 => std_logic_vector(to_unsigned( 128, 8)),
13 => std_logic_vector(to_unsigned( 70, 8)),
14 => std_logic_vector(to_unsigned( 80, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 22, 8)),
17 => std_logic_vector(to_unsigned( 52, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 924 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 4, 8)),
2 => std_logic_vector(to_unsigned( 184, 8)),
3 => std_logic_vector(to_unsigned( 195, 8)),
4 => std_logic_vector(to_unsigned( 253, 8)),
5 => std_logic_vector(to_unsigned( 145, 8)),
6 => std_logic_vector(to_unsigned( 57, 8)),
7 => std_logic_vector(to_unsigned( 26, 8)),
8 => std_logic_vector(to_unsigned( 167, 8)),
9 => std_logic_vector(to_unsigned( 162, 8)),
10 => std_logic_vector(to_unsigned( 40, 8)),
11 => std_logic_vector(to_unsigned( 146, 8)),
12 => std_logic_vector(to_unsigned( 56, 8)),
13 => std_logic_vector(to_unsigned( 249, 8)),
14 => std_logic_vector(to_unsigned( 96, 8)),
15 => std_logic_vector(to_unsigned( 196, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 180, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 925 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 108, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 69, 8)),
4 => std_logic_vector(to_unsigned( 147, 8)),
5 => std_logic_vector(to_unsigned( 235, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 46, 8)),
8 => std_logic_vector(to_unsigned( 124, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 20, 8)),
12 => std_logic_vector(to_unsigned( 98, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 19, 8)),
15 => std_logic_vector(to_unsigned( 76, 8)),
16 => std_logic_vector(to_unsigned( 142, 8)),
17 => std_logic_vector(to_unsigned( 70, 8)),
18 => std_logic_vector(to_unsigned( 79, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 926 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 68, 8)),
2 => std_logic_vector(to_unsigned( 85, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 123, 8)),
5 => std_logic_vector(to_unsigned( 182, 8)),
6 => std_logic_vector(to_unsigned( 97, 8)),
7 => std_logic_vector(to_unsigned( 105, 8)),
8 => std_logic_vector(to_unsigned( 48, 8)),
9 => std_logic_vector(to_unsigned( 1, 8)),
10 => std_logic_vector(to_unsigned( 146, 8)),
11 => std_logic_vector(to_unsigned( 17, 8)),
12 => std_logic_vector(to_unsigned( 24, 8)),
13 => std_logic_vector(to_unsigned( 94, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 191, 8)),
16 => std_logic_vector(to_unsigned( 18, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 927 then RAM <= (0 => "01101111",
1 => std_logic_vector(to_unsigned( 46, 8)),
2 => std_logic_vector(to_unsigned( 98, 8)),
3 => std_logic_vector(to_unsigned( 104, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 30, 8)),
6 => std_logic_vector(to_unsigned( 120, 8)),
7 => std_logic_vector(to_unsigned( 62, 8)),
8 => std_logic_vector(to_unsigned( 152, 8)),
9 => std_logic_vector(to_unsigned( 119, 8)),
10 => std_logic_vector(to_unsigned( 183, 8)),
11 => std_logic_vector(to_unsigned( 69, 8)),
12 => std_logic_vector(to_unsigned( 75, 8)),
13 => std_logic_vector(to_unsigned( 62, 8)),
14 => std_logic_vector(to_unsigned( 205, 8)),
15 => std_logic_vector(to_unsigned( 53, 8)),
16 => std_logic_vector(to_unsigned( 160, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101101
elsif count = 928 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 177, 8)),
2 => std_logic_vector(to_unsigned( 102, 8)),
3 => std_logic_vector(to_unsigned( 173, 8)),
4 => std_logic_vector(to_unsigned( 98, 8)),
5 => std_logic_vector(to_unsigned( 245, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 135, 8)),
8 => std_logic_vector(to_unsigned( 134, 8)),
9 => std_logic_vector(to_unsigned( 194, 8)),
10 => std_logic_vector(to_unsigned( 151, 8)),
11 => std_logic_vector(to_unsigned( 32, 8)),
12 => std_logic_vector(to_unsigned( 207, 8)),
13 => std_logic_vector(to_unsigned( 204, 8)),
14 => std_logic_vector(to_unsigned( 141, 8)),
15 => std_logic_vector(to_unsigned( 139, 8)),
16 => std_logic_vector(to_unsigned( 140, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 929 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 83, 8)),
4 => std_logic_vector(to_unsigned( 101, 8)),
5 => std_logic_vector(to_unsigned( 16, 8)),
6 => std_logic_vector(to_unsigned( 67, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 158, 8)),
9 => std_logic_vector(to_unsigned( 108, 8)),
10 => std_logic_vector(to_unsigned( 208, 8)),
11 => std_logic_vector(to_unsigned( 126, 8)),
12 => std_logic_vector(to_unsigned( 190, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 101, 8)),
15 => std_logic_vector(to_unsigned( 242, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 151, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 930 then RAM <= (0 => "11010111",
1 => std_logic_vector(to_unsigned( 140, 8)),
2 => std_logic_vector(to_unsigned( 167, 8)),
3 => std_logic_vector(to_unsigned( 137, 8)),
4 => std_logic_vector(to_unsigned( 164, 8)),
5 => std_logic_vector(to_unsigned( 103, 8)),
6 => std_logic_vector(to_unsigned( 124, 8)),
7 => std_logic_vector(to_unsigned( 47, 8)),
8 => std_logic_vector(to_unsigned( 195, 8)),
9 => std_logic_vector(to_unsigned( 175, 8)),
10 => std_logic_vector(to_unsigned( 172, 8)),
11 => std_logic_vector(to_unsigned( 151, 8)),
12 => std_logic_vector(to_unsigned( 4, 8)),
13 => std_logic_vector(to_unsigned( 120, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 216, 8)),
16 => std_logic_vector(to_unsigned( 131, 8)),
17 => std_logic_vector(to_unsigned( 160, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010111
elsif count = 931 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 124, 8)),
3 => std_logic_vector(to_unsigned( 138, 8)),
4 => std_logic_vector(to_unsigned( 63, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 93, 8)),
8 => std_logic_vector(to_unsigned( 138, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 170, 8)),
11 => std_logic_vector(to_unsigned( 20, 8)),
12 => std_logic_vector(to_unsigned( 230, 8)),
13 => std_logic_vector(to_unsigned( 90, 8)),
14 => std_logic_vector(to_unsigned( 18, 8)),
15 => std_logic_vector(to_unsigned( 123, 8)),
16 => std_logic_vector(to_unsigned( 168, 8)),
17 => std_logic_vector(to_unsigned( 153, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011110
elsif count = 932 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 194, 8)),
2 => std_logic_vector(to_unsigned( 154, 8)),
3 => std_logic_vector(to_unsigned( 148, 8)),
4 => std_logic_vector(to_unsigned( 82, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 237, 8)),
8 => std_logic_vector(to_unsigned( 163, 8)),
9 => std_logic_vector(to_unsigned( 189, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 202, 8)),
12 => std_logic_vector(to_unsigned( 94, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 128, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 155, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010001
elsif count = 933 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 13, 8)),
2 => std_logic_vector(to_unsigned( 56, 8)),
3 => std_logic_vector(to_unsigned( 24, 8)),
4 => std_logic_vector(to_unsigned( 105, 8)),
5 => std_logic_vector(to_unsigned( 98, 8)),
6 => std_logic_vector(to_unsigned( 175, 8)),
7 => std_logic_vector(to_unsigned( 131, 8)),
8 => std_logic_vector(to_unsigned( 142, 8)),
9 => std_logic_vector(to_unsigned( 254, 8)),
10 => std_logic_vector(to_unsigned( 236, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 61, 8)),
13 => std_logic_vector(to_unsigned( 203, 8)),
14 => std_logic_vector(to_unsigned( 53, 8)),
15 => std_logic_vector(to_unsigned( 160, 8)),
16 => std_logic_vector(to_unsigned( 113, 8)),
17 => std_logic_vector(to_unsigned( 96, 8)),
18 => std_logic_vector(to_unsigned( 102, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001110
elsif count = 934 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 115, 8)),
2 => std_logic_vector(to_unsigned( 84, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 124, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 88, 8)),
7 => std_logic_vector(to_unsigned( 82, 8)),
8 => std_logic_vector(to_unsigned( 157, 8)),
9 => std_logic_vector(to_unsigned( 228, 8)),
10 => std_logic_vector(to_unsigned( 49, 8)),
11 => std_logic_vector(to_unsigned( 175, 8)),
12 => std_logic_vector(to_unsigned( 150, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 227, 8)),
15 => std_logic_vector(to_unsigned( 101, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 113, 8)),
18 => std_logic_vector(to_unsigned( 135, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10001111
elsif count = 935 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 86, 8)),
2 => std_logic_vector(to_unsigned( 44, 8)),
3 => std_logic_vector(to_unsigned( 32, 8)),
4 => std_logic_vector(to_unsigned( 46, 8)),
5 => std_logic_vector(to_unsigned( 62, 8)),
6 => std_logic_vector(to_unsigned( 112, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 57, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 24, 8)),
12 => std_logic_vector(to_unsigned( 78, 8)),
13 => std_logic_vector(to_unsigned( 86, 8)),
14 => std_logic_vector(to_unsigned( 228, 8)),
15 => std_logic_vector(to_unsigned( 40, 8)),
16 => std_logic_vector(to_unsigned( 38, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 66, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 936 then RAM <= (0 => "10101111",
1 => std_logic_vector(to_unsigned( 143, 8)),
2 => std_logic_vector(to_unsigned( 130, 8)),
3 => std_logic_vector(to_unsigned( 196, 8)),
4 => std_logic_vector(to_unsigned( 35, 8)),
5 => std_logic_vector(to_unsigned( 108, 8)),
6 => std_logic_vector(to_unsigned( 75, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 69, 8)),
10 => std_logic_vector(to_unsigned( 24, 8)),
11 => std_logic_vector(to_unsigned( 232, 8)),
12 => std_logic_vector(to_unsigned( 99, 8)),
13 => std_logic_vector(to_unsigned( 94, 8)),
14 => std_logic_vector(to_unsigned( 176, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 104, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 937 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 153, 8)),
3 => std_logic_vector(to_unsigned( 93, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 39, 8)),
6 => std_logic_vector(to_unsigned( 140, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 104, 8)),
9 => std_logic_vector(to_unsigned( 196, 8)),
10 => std_logic_vector(to_unsigned( 161, 8)),
11 => std_logic_vector(to_unsigned( 232, 8)),
12 => std_logic_vector(to_unsigned( 65, 8)),
13 => std_logic_vector(to_unsigned( 91, 8)),
14 => std_logic_vector(to_unsigned( 140, 8)),
15 => std_logic_vector(to_unsigned( 240, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 65, 8)),
18 => std_logic_vector(to_unsigned( 104, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 938 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 7, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 36, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 74, 8)),
6 => std_logic_vector(to_unsigned( 142, 8)),
7 => std_logic_vector(to_unsigned( 40, 8)),
8 => std_logic_vector(to_unsigned( 108, 8)),
9 => std_logic_vector(to_unsigned( 28, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 27, 8)),
13 => std_logic_vector(to_unsigned( 56, 8)),
14 => std_logic_vector(to_unsigned( 124, 8)),
15 => std_logic_vector(to_unsigned( 85, 8)),
16 => std_logic_vector(to_unsigned( 33, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001100
elsif count = 939 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 224, 8)),
2 => std_logic_vector(to_unsigned( 195, 8)),
3 => std_logic_vector(to_unsigned( 105, 8)),
4 => std_logic_vector(to_unsigned( 17, 8)),
5 => std_logic_vector(to_unsigned( 31, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 200, 8)),
8 => std_logic_vector(to_unsigned( 178, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 65, 8)),
11 => std_logic_vector(to_unsigned( 54, 8)),
12 => std_logic_vector(to_unsigned( 54, 8)),
13 => std_logic_vector(to_unsigned( 75, 8)),
14 => std_logic_vector(to_unsigned( 109, 8)),
15 => std_logic_vector(to_unsigned( 73, 8)),
16 => std_logic_vector(to_unsigned( 35, 8)),
17 => std_logic_vector(to_unsigned( 98, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110010
elsif count = 940 then RAM <= (0 => "01111011",
1 => std_logic_vector(to_unsigned( 79, 8)),
2 => std_logic_vector(to_unsigned( 97, 8)),
3 => std_logic_vector(to_unsigned( 95, 8)),
4 => std_logic_vector(to_unsigned( 75, 8)),
5 => std_logic_vector(to_unsigned( 50, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 134, 8)),
8 => std_logic_vector(to_unsigned( 36, 8)),
9 => std_logic_vector(to_unsigned( 169, 8)),
10 => std_logic_vector(to_unsigned( 41, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 61, 8)),
13 => std_logic_vector(to_unsigned( 115, 8)),
14 => std_logic_vector(to_unsigned( 133, 8)),
15 => std_logic_vector(to_unsigned( 179, 8)),
16 => std_logic_vector(to_unsigned( 247, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 941 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 96, 8)),
2 => std_logic_vector(to_unsigned( 76, 8)),
3 => std_logic_vector(to_unsigned( 179, 8)),
4 => std_logic_vector(to_unsigned( 154, 8)),
5 => std_logic_vector(to_unsigned( 232, 8)),
6 => std_logic_vector(to_unsigned( 77, 8)),
7 => std_logic_vector(to_unsigned( 142, 8)),
8 => std_logic_vector(to_unsigned( 242, 8)),
9 => std_logic_vector(to_unsigned( 158, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 232, 8)),
12 => std_logic_vector(to_unsigned( 33, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 136, 8)),
16 => std_logic_vector(to_unsigned( 135, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 89, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010110
elsif count = 942 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 5, 8)),
2 => std_logic_vector(to_unsigned( 114, 8)),
3 => std_logic_vector(to_unsigned( 108, 8)),
4 => std_logic_vector(to_unsigned( 169, 8)),
5 => std_logic_vector(to_unsigned( 70, 8)),
6 => std_logic_vector(to_unsigned( 82, 8)),
7 => std_logic_vector(to_unsigned( 109, 8)),
8 => std_logic_vector(to_unsigned( 62, 8)),
9 => std_logic_vector(to_unsigned( 196, 8)),
10 => std_logic_vector(to_unsigned( 157, 8)),
11 => std_logic_vector(to_unsigned( 214, 8)),
12 => std_logic_vector(to_unsigned( 8, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 105, 8)),
15 => std_logic_vector(to_unsigned( 110, 8)),
16 => std_logic_vector(to_unsigned( 171, 8)),
17 => std_logic_vector(to_unsigned( 146, 8)),
18 => std_logic_vector(to_unsigned( 142, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11010010
elsif count = 943 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 249, 8)),
3 => std_logic_vector(to_unsigned( 250, 8)),
4 => std_logic_vector(to_unsigned( 90, 8)),
5 => std_logic_vector(to_unsigned( 176, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 99, 8)),
8 => std_logic_vector(to_unsigned( 27, 8)),
9 => std_logic_vector(to_unsigned( 208, 8)),
10 => std_logic_vector(to_unsigned( 132, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 43, 8)),
13 => std_logic_vector(to_unsigned( 194, 8)),
14 => std_logic_vector(to_unsigned( 184, 8)),
15 => std_logic_vector(to_unsigned( 243, 8)),
16 => std_logic_vector(to_unsigned( 163, 8)),
17 => std_logic_vector(to_unsigned( 194, 8)),
18 => std_logic_vector(to_unsigned( 90, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00110110
elsif count = 944 then RAM <= (0 => "11111001",
1 => std_logic_vector(to_unsigned( 123, 8)),
2 => std_logic_vector(to_unsigned( 169, 8)),
3 => std_logic_vector(to_unsigned( 199, 8)),
4 => std_logic_vector(to_unsigned( 38, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 108, 8)),
7 => std_logic_vector(to_unsigned( 74, 8)),
8 => std_logic_vector(to_unsigned( 233, 8)),
9 => std_logic_vector(to_unsigned( 177, 8)),
10 => std_logic_vector(to_unsigned( 199, 8)),
11 => std_logic_vector(to_unsigned( 102, 8)),
12 => std_logic_vector(to_unsigned( 148, 8)),
13 => std_logic_vector(to_unsigned( 146, 8)),
14 => std_logic_vector(to_unsigned( 192, 8)),
15 => std_logic_vector(to_unsigned( 165, 8)),
16 => std_logic_vector(to_unsigned( 211, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 144, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110001
elsif count = 945 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 243, 8)),
3 => std_logic_vector(to_unsigned( 42, 8)),
4 => std_logic_vector(to_unsigned( 248, 8)),
5 => std_logic_vector(to_unsigned( 188, 8)),
6 => std_logic_vector(to_unsigned( 152, 8)),
7 => std_logic_vector(to_unsigned( 28, 8)),
8 => std_logic_vector(to_unsigned( 121, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 202, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 141, 8)),
13 => std_logic_vector(to_unsigned( 89, 8)),
14 => std_logic_vector(to_unsigned( 195, 8)),
15 => std_logic_vector(to_unsigned( 190, 8)),
16 => std_logic_vector(to_unsigned( 204, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 179, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 946 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 173, 8)),
3 => std_logic_vector(to_unsigned( 151, 8)),
4 => std_logic_vector(to_unsigned( 60, 8)),
5 => std_logic_vector(to_unsigned( 132, 8)),
6 => std_logic_vector(to_unsigned( 79, 8)),
7 => std_logic_vector(to_unsigned( 127, 8)),
8 => std_logic_vector(to_unsigned( 84, 8)),
9 => std_logic_vector(to_unsigned( 31, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 183, 8)),
12 => std_logic_vector(to_unsigned( 182, 8)),
13 => std_logic_vector(to_unsigned( 196, 8)),
14 => std_logic_vector(to_unsigned( 189, 8)),
15 => std_logic_vector(to_unsigned( 221, 8)),
16 => std_logic_vector(to_unsigned( 23, 8)),
17 => std_logic_vector(to_unsigned( 165, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 947 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 110, 8)),
3 => std_logic_vector(to_unsigned( 156, 8)),
4 => std_logic_vector(to_unsigned( 128, 8)),
5 => std_logic_vector(to_unsigned( 146, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 130, 8)),
8 => std_logic_vector(to_unsigned( 154, 8)),
9 => std_logic_vector(to_unsigned( 196, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 49, 8)),
13 => std_logic_vector(to_unsigned( 101, 8)),
14 => std_logic_vector(to_unsigned( 129, 8)),
15 => std_logic_vector(to_unsigned( 255, 8)),
16 => std_logic_vector(to_unsigned( 249, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 93, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101011
elsif count = 948 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 97, 8)),
2 => std_logic_vector(to_unsigned( 238, 8)),
3 => std_logic_vector(to_unsigned( 118, 8)),
4 => std_logic_vector(to_unsigned( 135, 8)),
5 => std_logic_vector(to_unsigned( 84, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 38, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 82, 8)),
10 => std_logic_vector(to_unsigned( 9, 8)),
11 => std_logic_vector(to_unsigned( 209, 8)),
12 => std_logic_vector(to_unsigned( 125, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 72, 8)),
16 => std_logic_vector(to_unsigned( 233, 8)),
17 => std_logic_vector(to_unsigned( 87, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 949 then RAM <= (0 => "11101011",
1 => std_logic_vector(to_unsigned( 58, 8)),
2 => std_logic_vector(to_unsigned( 254, 8)),
3 => std_logic_vector(to_unsigned( 240, 8)),
4 => std_logic_vector(to_unsigned( 173, 8)),
5 => std_logic_vector(to_unsigned( 138, 8)),
6 => std_logic_vector(to_unsigned( 129, 8)),
7 => std_logic_vector(to_unsigned( 79, 8)),
8 => std_logic_vector(to_unsigned( 233, 8)),
9 => std_logic_vector(to_unsigned( 241, 8)),
10 => std_logic_vector(to_unsigned( 118, 8)),
11 => std_logic_vector(to_unsigned( 86, 8)),
12 => std_logic_vector(to_unsigned( 226, 8)),
13 => std_logic_vector(to_unsigned( 26, 8)),
14 => std_logic_vector(to_unsigned( 222, 8)),
15 => std_logic_vector(to_unsigned( 46, 8)),
16 => std_logic_vector(to_unsigned( 158, 8)),
17 => std_logic_vector(to_unsigned( 58, 8)),
18 => std_logic_vector(to_unsigned( 200, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101001
elsif count = 950 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 106, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 132, 8)),
4 => std_logic_vector(to_unsigned( 146, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 141, 8)),
7 => std_logic_vector(to_unsigned( 91, 8)),
8 => std_logic_vector(to_unsigned( 209, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 55, 8)),
11 => std_logic_vector(to_unsigned( 174, 8)),
12 => std_logic_vector(to_unsigned( 137, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 169, 8)),
15 => std_logic_vector(to_unsigned( 202, 8)),
16 => std_logic_vector(to_unsigned( 183, 8)),
17 => std_logic_vector(to_unsigned( 99, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001111
elsif count = 951 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 67, 8)),
2 => std_logic_vector(to_unsigned( 11, 8)),
3 => std_logic_vector(to_unsigned( 54, 8)),
4 => std_logic_vector(to_unsigned( 151, 8)),
5 => std_logic_vector(to_unsigned( 81, 8)),
6 => std_logic_vector(to_unsigned( 178, 8)),
7 => std_logic_vector(to_unsigned( 18, 8)),
8 => std_logic_vector(to_unsigned( 70, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 17, 8)),
11 => std_logic_vector(to_unsigned( 31, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 60, 8)),
14 => std_logic_vector(to_unsigned( 227, 8)),
15 => std_logic_vector(to_unsigned( 21, 8)),
16 => std_logic_vector(to_unsigned( 184, 8)),
17 => std_logic_vector(to_unsigned( 54, 8)),
18 => std_logic_vector(to_unsigned( 192, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 952 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 180, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 194, 8)),
6 => std_logic_vector(to_unsigned( 107, 8)),
7 => std_logic_vector(to_unsigned( 205, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 225, 8)),
11 => std_logic_vector(to_unsigned( 104, 8)),
12 => std_logic_vector(to_unsigned( 102, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 84, 8)),
15 => std_logic_vector(to_unsigned( 197, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 166, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001111
elsif count = 953 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 73, 8)),
2 => std_logic_vector(to_unsigned( 161, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 152, 8)),
7 => std_logic_vector(to_unsigned( 113, 8)),
8 => std_logic_vector(to_unsigned( 43, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 233, 8)),
11 => std_logic_vector(to_unsigned( 22, 8)),
12 => std_logic_vector(to_unsigned( 107, 8)),
13 => std_logic_vector(to_unsigned( 98, 8)),
14 => std_logic_vector(to_unsigned( 164, 8)),
15 => std_logic_vector(to_unsigned( 83, 8)),
16 => std_logic_vector(to_unsigned( 211, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 181, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 954 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 144, 8)),
2 => std_logic_vector(to_unsigned( 103, 8)),
3 => std_logic_vector(to_unsigned( 250, 8)),
4 => std_logic_vector(to_unsigned( 121, 8)),
5 => std_logic_vector(to_unsigned( 144, 8)),
6 => std_logic_vector(to_unsigned( 103, 8)),
7 => std_logic_vector(to_unsigned( 121, 8)),
8 => std_logic_vector(to_unsigned( 126, 8)),
9 => std_logic_vector(to_unsigned( 192, 8)),
10 => std_logic_vector(to_unsigned( 220, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 72, 8)),
13 => std_logic_vector(to_unsigned( 104, 8)),
14 => std_logic_vector(to_unsigned( 111, 8)),
15 => std_logic_vector(to_unsigned( 122, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 120, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 955 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 185, 8)),
2 => std_logic_vector(to_unsigned( 151, 8)),
3 => std_logic_vector(to_unsigned( 53, 8)),
4 => std_logic_vector(to_unsigned( 9, 8)),
5 => std_logic_vector(to_unsigned( 187, 8)),
6 => std_logic_vector(to_unsigned( 143, 8)),
7 => std_logic_vector(to_unsigned( 123, 8)),
8 => std_logic_vector(to_unsigned( 203, 8)),
9 => std_logic_vector(to_unsigned( 249, 8)),
10 => std_logic_vector(to_unsigned( 243, 8)),
11 => std_logic_vector(to_unsigned( 156, 8)),
12 => std_logic_vector(to_unsigned( 112, 8)),
13 => std_logic_vector(to_unsigned( 69, 8)),
14 => std_logic_vector(to_unsigned( 143, 8)),
15 => std_logic_vector(to_unsigned( 68, 8)),
16 => std_logic_vector(to_unsigned( 148, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 956 then RAM <= (0 => "11100111",
1 => std_logic_vector(to_unsigned( 162, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 141, 8)),
4 => std_logic_vector(to_unsigned( 207, 8)),
5 => std_logic_vector(to_unsigned( 226, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 133, 8)),
8 => std_logic_vector(to_unsigned( 25, 8)),
9 => std_logic_vector(to_unsigned( 38, 8)),
10 => std_logic_vector(to_unsigned( 53, 8)),
11 => std_logic_vector(to_unsigned( 140, 8)),
12 => std_logic_vector(to_unsigned( 245, 8)),
13 => std_logic_vector(to_unsigned( 54, 8)),
14 => std_logic_vector(to_unsigned( 134, 8)),
15 => std_logic_vector(to_unsigned( 48, 8)),
16 => std_logic_vector(to_unsigned( 152, 8)),
17 => std_logic_vector(to_unsigned( 122, 8)),
18 => std_logic_vector(to_unsigned( 146, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11000011
elsif count = 957 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 111, 8)),
2 => std_logic_vector(to_unsigned( 65, 8)),
3 => std_logic_vector(to_unsigned( 83, 8)),
4 => std_logic_vector(to_unsigned( 99, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 215, 8)),
7 => std_logic_vector(to_unsigned( 96, 8)),
8 => std_logic_vector(to_unsigned( 50, 8)),
9 => std_logic_vector(to_unsigned( 122, 8)),
10 => std_logic_vector(to_unsigned( 50, 8)),
11 => std_logic_vector(to_unsigned( 55, 8)),
12 => std_logic_vector(to_unsigned( 71, 8)),
13 => std_logic_vector(to_unsigned( 61, 8)),
14 => std_logic_vector(to_unsigned( 77, 8)),
15 => std_logic_vector(to_unsigned( 112, 8)),
16 => std_logic_vector(to_unsigned( 66, 8)),
17 => std_logic_vector(to_unsigned( 83, 8)),
18 => std_logic_vector(to_unsigned( 68, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101011
elsif count = 958 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 66, 8)),
2 => std_logic_vector(to_unsigned( 232, 8)),
3 => std_logic_vector(to_unsigned( 189, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 253, 8)),
6 => std_logic_vector(to_unsigned( 214, 8)),
7 => std_logic_vector(to_unsigned( 181, 8)),
8 => std_logic_vector(to_unsigned( 212, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 211, 8)),
13 => std_logic_vector(to_unsigned( 204, 8)),
14 => std_logic_vector(to_unsigned( 27, 8)),
15 => std_logic_vector(to_unsigned( 133, 8)),
16 => std_logic_vector(to_unsigned( 117, 8)),
17 => std_logic_vector(to_unsigned( 171, 8)),
18 => std_logic_vector(to_unsigned( 176, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111010
elsif count = 959 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 223, 8)),
2 => std_logic_vector(to_unsigned( 44, 8)),
3 => std_logic_vector(to_unsigned( 116, 8)),
4 => std_logic_vector(to_unsigned( 136, 8)),
5 => std_logic_vector(to_unsigned( 125, 8)),
6 => std_logic_vector(to_unsigned( 145, 8)),
7 => std_logic_vector(to_unsigned( 125, 8)),
8 => std_logic_vector(to_unsigned( 79, 8)),
9 => std_logic_vector(to_unsigned( 209, 8)),
10 => std_logic_vector(to_unsigned( 149, 8)),
11 => std_logic_vector(to_unsigned( 118, 8)),
12 => std_logic_vector(to_unsigned( 86, 8)),
13 => std_logic_vector(to_unsigned( 6, 8)),
14 => std_logic_vector(to_unsigned( 43, 8)),
15 => std_logic_vector(to_unsigned( 95, 8)),
16 => std_logic_vector(to_unsigned( 109, 8)),
17 => std_logic_vector(to_unsigned( 169, 8)),
18 => std_logic_vector(to_unsigned( 112, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10111110
elsif count = 960 then RAM <= (0 => "11111110",
1 => std_logic_vector(to_unsigned( 154, 8)),
2 => std_logic_vector(to_unsigned( 234, 8)),
3 => std_logic_vector(to_unsigned( 113, 8)),
4 => std_logic_vector(to_unsigned( 99, 8)),
5 => std_logic_vector(to_unsigned( 181, 8)),
6 => std_logic_vector(to_unsigned( 138, 8)),
7 => std_logic_vector(to_unsigned( 154, 8)),
8 => std_logic_vector(to_unsigned( 58, 8)),
9 => std_logic_vector(to_unsigned( 129, 8)),
10 => std_logic_vector(to_unsigned( 21, 8)),
11 => std_logic_vector(to_unsigned( 84, 8)),
12 => std_logic_vector(to_unsigned( 0, 8)),
13 => std_logic_vector(to_unsigned( 85, 8)),
14 => std_logic_vector(to_unsigned( 79, 8)),
15 => std_logic_vector(to_unsigned( 75, 8)),
16 => std_logic_vector(to_unsigned( 69, 8)),
17 => std_logic_vector(to_unsigned( 109, 8)),
18 => std_logic_vector(to_unsigned( 52, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 961 then RAM <= (0 => "11001111",
1 => std_logic_vector(to_unsigned( 126, 8)),
2 => std_logic_vector(to_unsigned( 106, 8)),
3 => std_logic_vector(to_unsigned( 149, 8)),
4 => std_logic_vector(to_unsigned( 109, 8)),
5 => std_logic_vector(to_unsigned( 195, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 119, 8)),
8 => std_logic_vector(to_unsigned( 113, 8)),
9 => std_logic_vector(to_unsigned( 207, 8)),
10 => std_logic_vector(to_unsigned( 169, 8)),
11 => std_logic_vector(to_unsigned( 78, 8)),
12 => std_logic_vector(to_unsigned( 12, 8)),
13 => std_logic_vector(to_unsigned( 143, 8)),
14 => std_logic_vector(to_unsigned( 173, 8)),
15 => std_logic_vector(to_unsigned( 201, 8)),
16 => std_logic_vector(to_unsigned( 67, 8)),
17 => std_logic_vector(to_unsigned( 136, 8)),
18 => std_logic_vector(to_unsigned( 138, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01001011
elsif count = 962 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 155, 8)),
2 => std_logic_vector(to_unsigned( 88, 8)),
3 => std_logic_vector(to_unsigned( 135, 8)),
4 => std_logic_vector(to_unsigned( 108, 8)),
5 => std_logic_vector(to_unsigned( 160, 8)),
6 => std_logic_vector(to_unsigned( 205, 8)),
7 => std_logic_vector(to_unsigned( 182, 8)),
8 => std_logic_vector(to_unsigned( 81, 8)),
9 => std_logic_vector(to_unsigned( 42, 8)),
10 => std_logic_vector(to_unsigned( 42, 8)),
11 => std_logic_vector(to_unsigned( 143, 8)),
12 => std_logic_vector(to_unsigned( 118, 8)),
13 => std_logic_vector(to_unsigned( 131, 8)),
14 => std_logic_vector(to_unsigned( 198, 8)),
15 => std_logic_vector(to_unsigned( 22, 8)),
16 => std_logic_vector(to_unsigned( 234, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 109, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101011
elsif count = 963 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 38, 8)),
2 => std_logic_vector(to_unsigned( 66, 8)),
3 => std_logic_vector(to_unsigned( 88, 8)),
4 => std_logic_vector(to_unsigned( 38, 8)),
5 => std_logic_vector(to_unsigned( 36, 8)),
6 => std_logic_vector(to_unsigned( 64, 8)),
7 => std_logic_vector(to_unsigned( 252, 8)),
8 => std_logic_vector(to_unsigned( 97, 8)),
9 => std_logic_vector(to_unsigned( 64, 8)),
10 => std_logic_vector(to_unsigned( 14, 8)),
11 => std_logic_vector(to_unsigned( 66, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 88, 8)),
14 => std_logic_vector(to_unsigned( 38, 8)),
15 => std_logic_vector(to_unsigned( 212, 8)),
16 => std_logic_vector(to_unsigned( 224, 8)),
17 => std_logic_vector(to_unsigned( 60, 8)),
18 => std_logic_vector(to_unsigned( 49, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110111
elsif count = 964 then RAM <= (0 => "11101110",
1 => std_logic_vector(to_unsigned( 121, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 125, 8)),
4 => std_logic_vector(to_unsigned( 122, 8)),
5 => std_logic_vector(to_unsigned( 69, 8)),
6 => std_logic_vector(to_unsigned( 162, 8)),
7 => std_logic_vector(to_unsigned( 204, 8)),
8 => std_logic_vector(to_unsigned( 236, 8)),
9 => std_logic_vector(to_unsigned( 22, 8)),
10 => std_logic_vector(to_unsigned( 152, 8)),
11 => std_logic_vector(to_unsigned( 47, 8)),
12 => std_logic_vector(to_unsigned( 140, 8)),
13 => std_logic_vector(to_unsigned( 99, 8)),
14 => std_logic_vector(to_unsigned( 148, 8)),
15 => std_logic_vector(to_unsigned( 72, 8)),
16 => std_logic_vector(to_unsigned( 165, 8)),
17 => std_logic_vector(to_unsigned( 77, 8)),
18 => std_logic_vector(to_unsigned( 117, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100110
elsif count = 965 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 193, 8)),
2 => std_logic_vector(to_unsigned( 237, 8)),
3 => std_logic_vector(to_unsigned( 162, 8)),
4 => std_logic_vector(to_unsigned( 208, 8)),
5 => std_logic_vector(to_unsigned( 154, 8)),
6 => std_logic_vector(to_unsigned( 85, 8)),
7 => std_logic_vector(to_unsigned( 162, 8)),
8 => std_logic_vector(to_unsigned( 208, 8)),
9 => std_logic_vector(to_unsigned( 150, 8)),
10 => std_logic_vector(to_unsigned( 230, 8)),
11 => std_logic_vector(to_unsigned( 122, 8)),
12 => std_logic_vector(to_unsigned( 120, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 223, 8)),
15 => std_logic_vector(to_unsigned( 28, 8)),
16 => std_logic_vector(to_unsigned( 79, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 225, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01011011
elsif count = 966 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 151, 8)),
2 => std_logic_vector(to_unsigned( 142, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 138, 8)),
5 => std_logic_vector(to_unsigned( 210, 8)),
6 => std_logic_vector(to_unsigned( 81, 8)),
7 => std_logic_vector(to_unsigned( 129, 8)),
8 => std_logic_vector(to_unsigned( 120, 8)),
9 => std_logic_vector(to_unsigned( 125, 8)),
10 => std_logic_vector(to_unsigned( 72, 8)),
11 => std_logic_vector(to_unsigned( 169, 8)),
12 => std_logic_vector(to_unsigned( 53, 8)),
13 => std_logic_vector(to_unsigned( 130, 8)),
14 => std_logic_vector(to_unsigned( 121, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 115, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 967 then RAM <= (0 => "01111101",
1 => std_logic_vector(to_unsigned( 146, 8)),
2 => std_logic_vector(to_unsigned( 100, 8)),
3 => std_logic_vector(to_unsigned( 16, 8)),
4 => std_logic_vector(to_unsigned( 186, 8)),
5 => std_logic_vector(to_unsigned( 136, 8)),
6 => std_logic_vector(to_unsigned( 110, 8)),
7 => std_logic_vector(to_unsigned( 68, 8)),
8 => std_logic_vector(to_unsigned( 54, 8)),
9 => std_logic_vector(to_unsigned( 32, 8)),
10 => std_logic_vector(to_unsigned( 110, 8)),
11 => std_logic_vector(to_unsigned( 136, 8)),
12 => std_logic_vector(to_unsigned( 90, 8)),
13 => std_logic_vector(to_unsigned( 145, 8)),
14 => std_logic_vector(to_unsigned( 99, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 139, 8)),
17 => std_logic_vector(to_unsigned( 84, 8)),
18 => std_logic_vector(to_unsigned( 100, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111101
elsif count = 968 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 114, 8)),
2 => std_logic_vector(to_unsigned( 61, 8)),
3 => std_logic_vector(to_unsigned( 193, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 111, 8)),
6 => std_logic_vector(to_unsigned( 218, 8)),
7 => std_logic_vector(to_unsigned( 115, 8)),
8 => std_logic_vector(to_unsigned( 220, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 60, 8)),
11 => std_logic_vector(to_unsigned( 76, 8)),
12 => std_logic_vector(to_unsigned( 183, 8)),
13 => std_logic_vector(to_unsigned( 103, 8)),
14 => std_logic_vector(to_unsigned( 210, 8)),
15 => std_logic_vector(to_unsigned( 182, 8)),
16 => std_logic_vector(to_unsigned( 129, 8)),
17 => std_logic_vector(to_unsigned( 114, 8)),
18 => std_logic_vector(to_unsigned( 141, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 969 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 159, 8)),
2 => std_logic_vector(to_unsigned( 95, 8)),
3 => std_logic_vector(to_unsigned( 130, 8)),
4 => std_logic_vector(to_unsigned( 43, 8)),
5 => std_logic_vector(to_unsigned( 181, 8)),
6 => std_logic_vector(to_unsigned( 139, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 252, 8)),
9 => std_logic_vector(to_unsigned( 25, 8)),
10 => std_logic_vector(to_unsigned( 253, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 117, 8)),
13 => std_logic_vector(to_unsigned( 229, 8)),
14 => std_logic_vector(to_unsigned( 40, 8)),
15 => std_logic_vector(to_unsigned( 186, 8)),
16 => std_logic_vector(to_unsigned( 122, 8)),
17 => std_logic_vector(to_unsigned( 129, 8)),
18 => std_logic_vector(to_unsigned( 128, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100101
elsif count = 970 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 188, 8)),
3 => std_logic_vector(to_unsigned( 71, 8)),
4 => std_logic_vector(to_unsigned( 198, 8)),
5 => std_logic_vector(to_unsigned( 54, 8)),
6 => std_logic_vector(to_unsigned( 240, 8)),
7 => std_logic_vector(to_unsigned( 118, 8)),
8 => std_logic_vector(to_unsigned( 199, 8)),
9 => std_logic_vector(to_unsigned( 71, 8)),
10 => std_logic_vector(to_unsigned( 198, 8)),
11 => std_logic_vector(to_unsigned( 89, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 107, 8)),
14 => std_logic_vector(to_unsigned( 170, 8)),
15 => std_logic_vector(to_unsigned( 37, 8)),
16 => std_logic_vector(to_unsigned( 72, 8)),
17 => std_logic_vector(to_unsigned( 95, 8)),
18 => std_logic_vector(to_unsigned( 190, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01111011
elsif count = 971 then RAM <= (0 => "10111111",
1 => std_logic_vector(to_unsigned( 93, 8)),
2 => std_logic_vector(to_unsigned( 108, 8)),
3 => std_logic_vector(to_unsigned( 115, 8)),
4 => std_logic_vector(to_unsigned( 114, 8)),
5 => std_logic_vector(to_unsigned( 92, 8)),
6 => std_logic_vector(to_unsigned( 237, 8)),
7 => std_logic_vector(to_unsigned( 90, 8)),
8 => std_logic_vector(to_unsigned( 111, 8)),
9 => std_logic_vector(to_unsigned( 193, 8)),
10 => std_logic_vector(to_unsigned( 124, 8)),
11 => std_logic_vector(to_unsigned( 162, 8)),
12 => std_logic_vector(to_unsigned( 161, 8)),
13 => std_logic_vector(to_unsigned( 149, 8)),
14 => std_logic_vector(to_unsigned( 127, 8)),
15 => std_logic_vector(to_unsigned( 92, 8)),
16 => std_logic_vector(to_unsigned( 237, 8)),
17 => std_logic_vector(to_unsigned( 101, 8)),
18 => std_logic_vector(to_unsigned( 173, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101111
elsif count = 972 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 172, 8)),
3 => std_logic_vector(to_unsigned( 52, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 140, 8)),
6 => std_logic_vector(to_unsigned( 181, 8)),
7 => std_logic_vector(to_unsigned( 117, 8)),
8 => std_logic_vector(to_unsigned( 204, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 194, 8)),
11 => std_logic_vector(to_unsigned( 117, 8)),
12 => std_logic_vector(to_unsigned( 119, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 70, 8)),
15 => std_logic_vector(to_unsigned( 217, 8)),
16 => std_logic_vector(to_unsigned( 105, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 165, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011111
elsif count = 973 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 149, 8)),
2 => std_logic_vector(to_unsigned( 210, 8)),
3 => std_logic_vector(to_unsigned( 203, 8)),
4 => std_logic_vector(to_unsigned( 123, 8)),
5 => std_logic_vector(to_unsigned( 107, 8)),
6 => std_logic_vector(to_unsigned( 35, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 140, 8)),
9 => std_logic_vector(to_unsigned( 20, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 177, 8)),
12 => std_logic_vector(to_unsigned( 61, 8)),
13 => std_logic_vector(to_unsigned( 125, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 72, 8)),
16 => std_logic_vector(to_unsigned( 82, 8)),
17 => std_logic_vector(to_unsigned( 172, 8)),
18 => std_logic_vector(to_unsigned( 105, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01101010
elsif count = 974 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 35, 8)),
2 => std_logic_vector(to_unsigned( 207, 8)),
3 => std_logic_vector(to_unsigned( 22, 8)),
4 => std_logic_vector(to_unsigned( 59, 8)),
5 => std_logic_vector(to_unsigned( 85, 8)),
6 => std_logic_vector(to_unsigned( 155, 8)),
7 => std_logic_vector(to_unsigned( 120, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 206, 8)),
10 => std_logic_vector(to_unsigned( 181, 8)),
11 => std_logic_vector(to_unsigned( 61, 8)),
12 => std_logic_vector(to_unsigned( 174, 8)),
13 => std_logic_vector(to_unsigned( 93, 8)),
14 => std_logic_vector(to_unsigned( 163, 8)),
15 => std_logic_vector(to_unsigned( 158, 8)),
16 => std_logic_vector(to_unsigned( 110, 8)),
17 => std_logic_vector(to_unsigned( 141, 8)),
18 => std_logic_vector(to_unsigned( 152, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001100
elsif count = 975 then RAM <= (0 => "01111111",
1 => std_logic_vector(to_unsigned( 109, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 121, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 174, 8)),
6 => std_logic_vector(to_unsigned( 52, 8)),
7 => std_logic_vector(to_unsigned( 168, 8)),
8 => std_logic_vector(to_unsigned( 96, 8)),
9 => std_logic_vector(to_unsigned( 213, 8)),
10 => std_logic_vector(to_unsigned( 204, 8)),
11 => std_logic_vector(to_unsigned( 185, 8)),
12 => std_logic_vector(to_unsigned( 63, 8)),
13 => std_logic_vector(to_unsigned( 17, 8)),
14 => std_logic_vector(to_unsigned( 74, 8)),
15 => std_logic_vector(to_unsigned( 18, 8)),
16 => std_logic_vector(to_unsigned( 147, 8)),
17 => std_logic_vector(to_unsigned( 137, 8)),
18 => std_logic_vector(to_unsigned( 71, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00101111
elsif count = 976 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 51, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 230, 8)),
4 => std_logic_vector(to_unsigned( 115, 8)),
5 => std_logic_vector(to_unsigned( 9, 8)),
6 => std_logic_vector(to_unsigned( 41, 8)),
7 => std_logic_vector(to_unsigned( 157, 8)),
8 => std_logic_vector(to_unsigned( 176, 8)),
9 => std_logic_vector(to_unsigned( 211, 8)),
10 => std_logic_vector(to_unsigned( 93, 8)),
11 => std_logic_vector(to_unsigned( 20, 8)),
12 => std_logic_vector(to_unsigned( 152, 8)),
13 => std_logic_vector(to_unsigned( 139, 8)),
14 => std_logic_vector(to_unsigned( 158, 8)),
15 => std_logic_vector(to_unsigned( 123, 8)),
16 => std_logic_vector(to_unsigned( 112, 8)),
17 => std_logic_vector(to_unsigned( 175, 8)),
18 => std_logic_vector(to_unsigned( 127, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001010
elsif count = 977 then RAM <= (0 => "10011111",
1 => std_logic_vector(to_unsigned( 137, 8)),
2 => std_logic_vector(to_unsigned( 43, 8)),
3 => std_logic_vector(to_unsigned( 97, 8)),
4 => std_logic_vector(to_unsigned( 83, 8)),
5 => std_logic_vector(to_unsigned( 128, 8)),
6 => std_logic_vector(to_unsigned( 116, 8)),
7 => std_logic_vector(to_unsigned( 138, 8)),
8 => std_logic_vector(to_unsigned( 42, 8)),
9 => std_logic_vector(to_unsigned( 180, 8)),
10 => std_logic_vector(to_unsigned( 14, 8)),
11 => std_logic_vector(to_unsigned( 25, 8)),
12 => std_logic_vector(to_unsigned( 82, 8)),
13 => std_logic_vector(to_unsigned( 117, 8)),
14 => std_logic_vector(to_unsigned( 55, 8)),
15 => std_logic_vector(to_unsigned( 120, 8)),
16 => std_logic_vector(to_unsigned( 60, 8)),
17 => std_logic_vector(to_unsigned( 173, 8)),
18 => std_logic_vector(to_unsigned( 84, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10011111
elsif count = 978 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 212, 8)),
2 => std_logic_vector(to_unsigned( 3, 8)),
3 => std_logic_vector(to_unsigned( 68, 8)),
4 => std_logic_vector(to_unsigned( 31, 8)),
5 => std_logic_vector(to_unsigned( 117, 8)),
6 => std_logic_vector(to_unsigned( 163, 8)),
7 => std_logic_vector(to_unsigned( 225, 8)),
8 => std_logic_vector(to_unsigned( 168, 8)),
9 => std_logic_vector(to_unsigned( 27, 8)),
10 => std_logic_vector(to_unsigned( 14, 8)),
11 => std_logic_vector(to_unsigned( 9, 8)),
12 => std_logic_vector(to_unsigned( 32, 8)),
13 => std_logic_vector(to_unsigned( 53, 8)),
14 => std_logic_vector(to_unsigned( 16, 8)),
15 => std_logic_vector(to_unsigned( 174, 8)),
16 => std_logic_vector(to_unsigned( 120, 8)),
17 => std_logic_vector(to_unsigned( 39, 8)),
18 => std_logic_vector(to_unsigned( 40, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
elsif count = 979 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 153, 8)),
2 => std_logic_vector(to_unsigned( 174, 8)),
3 => std_logic_vector(to_unsigned( 74, 8)),
4 => std_logic_vector(to_unsigned( 224, 8)),
5 => std_logic_vector(to_unsigned( 45, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 87, 8)),
8 => std_logic_vector(to_unsigned( 116, 8)),
9 => std_logic_vector(to_unsigned( 146, 8)),
10 => std_logic_vector(to_unsigned( 175, 8)),
11 => std_logic_vector(to_unsigned( 182, 8)),
12 => std_logic_vector(to_unsigned( 51, 8)),
13 => std_logic_vector(to_unsigned( 13, 8)),
14 => std_logic_vector(to_unsigned( 60, 8)),
15 => std_logic_vector(to_unsigned( 111, 8)),
16 => std_logic_vector(to_unsigned( 45, 8)),
17 => std_logic_vector(to_unsigned( 149, 8)),
18 => std_logic_vector(to_unsigned( 98, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111001
elsif count = 980 then RAM <= (0 => "11101111",
1 => std_logic_vector(to_unsigned( 78, 8)),
2 => std_logic_vector(to_unsigned( 223, 8)),
3 => std_logic_vector(to_unsigned( 225, 8)),
4 => std_logic_vector(to_unsigned( 222, 8)),
5 => std_logic_vector(to_unsigned( 37, 8)),
6 => std_logic_vector(to_unsigned( 184, 8)),
7 => std_logic_vector(to_unsigned( 54, 8)),
8 => std_logic_vector(to_unsigned( 247, 8)),
9 => std_logic_vector(to_unsigned( 46, 8)),
10 => std_logic_vector(to_unsigned( 46, 8)),
11 => std_logic_vector(to_unsigned( 145, 8)),
12 => std_logic_vector(to_unsigned( 149, 8)),
13 => std_logic_vector(to_unsigned( 13, 8)),
14 => std_logic_vector(to_unsigned( 208, 8)),
15 => std_logic_vector(to_unsigned( 29, 8)),
16 => std_logic_vector(to_unsigned( 192, 8)),
17 => std_logic_vector(to_unsigned( 46, 8)),
18 => std_logic_vector(to_unsigned( 215, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 981 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 100, 8)),
2 => std_logic_vector(to_unsigned( 182, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 180, 8)),
5 => std_logic_vector(to_unsigned( 104, 8)),
6 => std_logic_vector(to_unsigned( 180, 8)),
7 => std_logic_vector(to_unsigned( 132, 8)),
8 => std_logic_vector(to_unsigned( 87, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 191, 8)),
11 => std_logic_vector(to_unsigned( 222, 8)),
12 => std_logic_vector(to_unsigned( 27, 8)),
13 => std_logic_vector(to_unsigned( 105, 8)),
14 => std_logic_vector(to_unsigned( 4, 8)),
15 => std_logic_vector(to_unsigned( 251, 8)),
16 => std_logic_vector(to_unsigned( 195, 8)),
17 => std_logic_vector(to_unsigned( 103, 8)),
18 => std_logic_vector(to_unsigned( 210, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00010111
elsif count = 982 then RAM <= (0 => "10111110",
1 => std_logic_vector(to_unsigned( 2, 8)),
2 => std_logic_vector(to_unsigned( 168, 8)),
3 => std_logic_vector(to_unsigned( 182, 8)),
4 => std_logic_vector(to_unsigned( 153, 8)),
5 => std_logic_vector(to_unsigned( 135, 8)),
6 => std_logic_vector(to_unsigned( 136, 8)),
7 => std_logic_vector(to_unsigned( 149, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 153, 8)),
10 => std_logic_vector(to_unsigned( 112, 8)),
11 => std_logic_vector(to_unsigned( 85, 8)),
12 => std_logic_vector(to_unsigned( 106, 8)),
13 => std_logic_vector(to_unsigned( 109, 8)),
14 => std_logic_vector(to_unsigned( 224, 8)),
15 => std_logic_vector(to_unsigned( 117, 8)),
16 => std_logic_vector(to_unsigned( 106, 8)),
17 => std_logic_vector(to_unsigned( 167, 8)),
18 => std_logic_vector(to_unsigned( 133, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00011110
elsif count = 983 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 57, 8)),
3 => std_logic_vector(to_unsigned( 216, 8)),
4 => std_logic_vector(to_unsigned( 163, 8)),
5 => std_logic_vector(to_unsigned( 155, 8)),
6 => std_logic_vector(to_unsigned( 42, 8)),
7 => std_logic_vector(to_unsigned( 32, 8)),
8 => std_logic_vector(to_unsigned( 30, 8)),
9 => std_logic_vector(to_unsigned( 118, 8)),
10 => std_logic_vector(to_unsigned( 112, 8)),
11 => std_logic_vector(to_unsigned( 194, 8)),
12 => std_logic_vector(to_unsigned( 89, 8)),
13 => std_logic_vector(to_unsigned( 191, 8)),
14 => std_logic_vector(to_unsigned( 92, 8)),
15 => std_logic_vector(to_unsigned( 142, 8)),
16 => std_logic_vector(to_unsigned( 53, 8)),
17 => std_logic_vector(to_unsigned( 154, 8)),
18 => std_logic_vector(to_unsigned( 85, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100101
elsif count = 984 then RAM <= (0 => "11111010",
1 => std_logic_vector(to_unsigned( 224, 8)),
2 => std_logic_vector(to_unsigned( 213, 8)),
3 => std_logic_vector(to_unsigned( 25, 8)),
4 => std_logic_vector(to_unsigned( 158, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 102, 8)),
7 => std_logic_vector(to_unsigned( 29, 8)),
8 => std_logic_vector(to_unsigned( 162, 8)),
9 => std_logic_vector(to_unsigned( 234, 8)),
10 => std_logic_vector(to_unsigned( 22, 8)),
11 => std_logic_vector(to_unsigned( 113, 8)),
12 => std_logic_vector(to_unsigned( 164, 8)),
13 => std_logic_vector(to_unsigned( 174, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 79, 8)),
16 => std_logic_vector(to_unsigned( 102, 8)),
17 => std_logic_vector(to_unsigned( 72, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10101010
elsif count = 985 then RAM <= (0 => "11101101",
1 => std_logic_vector(to_unsigned( 175, 8)),
2 => std_logic_vector(to_unsigned( 107, 8)),
3 => std_logic_vector(to_unsigned( 60, 8)),
4 => std_logic_vector(to_unsigned( 225, 8)),
5 => std_logic_vector(to_unsigned( 162, 8)),
6 => std_logic_vector(to_unsigned( 94, 8)),
7 => std_logic_vector(to_unsigned( 185, 8)),
8 => std_logic_vector(to_unsigned( 117, 8)),
9 => std_logic_vector(to_unsigned( 91, 8)),
10 => std_logic_vector(to_unsigned( 102, 8)),
11 => std_logic_vector(to_unsigned( 155, 8)),
12 => std_logic_vector(to_unsigned( 87, 8)),
13 => std_logic_vector(to_unsigned( 193, 8)),
14 => std_logic_vector(to_unsigned( 125, 8)),
15 => std_logic_vector(to_unsigned( 134, 8)),
16 => std_logic_vector(to_unsigned( 94, 8)),
17 => std_logic_vector(to_unsigned( 148, 8)),
18 => std_logic_vector(to_unsigned( 131, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101101
elsif count = 986 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 219, 8)),
2 => std_logic_vector(to_unsigned( 120, 8)),
3 => std_logic_vector(to_unsigned( 94, 8)),
4 => std_logic_vector(to_unsigned( 38, 8)),
5 => std_logic_vector(to_unsigned( 121, 8)),
6 => std_logic_vector(to_unsigned( 70, 8)),
7 => std_logic_vector(to_unsigned( 202, 8)),
8 => std_logic_vector(to_unsigned( 183, 8)),
9 => std_logic_vector(to_unsigned( 111, 8)),
10 => std_logic_vector(to_unsigned( 80, 8)),
11 => std_logic_vector(to_unsigned( 70, 8)),
12 => std_logic_vector(to_unsigned( 30, 8)),
13 => std_logic_vector(to_unsigned( 172, 8)),
14 => std_logic_vector(to_unsigned( 167, 8)),
15 => std_logic_vector(to_unsigned( 161, 8)),
16 => std_logic_vector(to_unsigned( 236, 8)),
17 => std_logic_vector(to_unsigned( 157, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010101
elsif count = 987 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 189, 8)),
2 => std_logic_vector(to_unsigned( 179, 8)),
3 => std_logic_vector(to_unsigned( 199, 8)),
4 => std_logic_vector(to_unsigned( 93, 8)),
5 => std_logic_vector(to_unsigned( 234, 8)),
6 => std_logic_vector(to_unsigned( 146, 8)),
7 => std_logic_vector(to_unsigned( 116, 8)),
8 => std_logic_vector(to_unsigned( 229, 8)),
9 => std_logic_vector(to_unsigned( 227, 8)),
10 => std_logic_vector(to_unsigned( 153, 8)),
11 => std_logic_vector(to_unsigned( 187, 8)),
12 => std_logic_vector(to_unsigned( 97, 8)),
13 => std_logic_vector(to_unsigned( 168, 8)),
14 => std_logic_vector(to_unsigned( 36, 8)),
15 => std_logic_vector(to_unsigned( 214, 8)),
16 => std_logic_vector(to_unsigned( 166, 8)),
17 => std_logic_vector(to_unsigned( 195, 8)),
18 => std_logic_vector(to_unsigned( 137, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110111
elsif count = 988 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 125, 8)),
2 => std_logic_vector(to_unsigned( 246, 8)),
3 => std_logic_vector(to_unsigned( 139, 8)),
4 => std_logic_vector(to_unsigned( 86, 8)),
5 => std_logic_vector(to_unsigned( 56, 8)),
6 => std_logic_vector(to_unsigned( 86, 8)),
7 => std_logic_vector(to_unsigned( 167, 8)),
8 => std_logic_vector(to_unsigned( 114, 8)),
9 => std_logic_vector(to_unsigned( 134, 8)),
10 => std_logic_vector(to_unsigned( 81, 8)),
11 => std_logic_vector(to_unsigned( 62, 8)),
12 => std_logic_vector(to_unsigned( 159, 8)),
13 => std_logic_vector(to_unsigned( 110, 8)),
14 => std_logic_vector(to_unsigned( 207, 8)),
15 => std_logic_vector(to_unsigned( 116, 8)),
16 => std_logic_vector(to_unsigned( 87, 8)),
17 => std_logic_vector(to_unsigned( 128, 8)),
18 => std_logic_vector(to_unsigned( 150, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11111010
elsif count = 989 then RAM <= (0 => "11011111",
1 => std_logic_vector(to_unsigned( 234, 8)),
2 => std_logic_vector(to_unsigned( 6, 8)),
3 => std_logic_vector(to_unsigned( 187, 8)),
4 => std_logic_vector(to_unsigned( 26, 8)),
5 => std_logic_vector(to_unsigned( 230, 8)),
6 => std_logic_vector(to_unsigned( 69, 8)),
7 => std_logic_vector(to_unsigned( 89, 8)),
8 => std_logic_vector(to_unsigned( 92, 8)),
9 => std_logic_vector(to_unsigned( 127, 8)),
10 => std_logic_vector(to_unsigned( 112, 8)),
11 => std_logic_vector(to_unsigned( 97, 8)),
12 => std_logic_vector(to_unsigned( 81, 8)),
13 => std_logic_vector(to_unsigned( 206, 8)),
14 => std_logic_vector(to_unsigned( 45, 8)),
15 => std_logic_vector(to_unsigned( 126, 8)),
16 => std_logic_vector(to_unsigned( 47, 8)),
17 => std_logic_vector(to_unsigned( 182, 8)),
18 => std_logic_vector(to_unsigned( 94, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01010110
elsif count = 990 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 41, 8)),
2 => std_logic_vector(to_unsigned( 19, 8)),
3 => std_logic_vector(to_unsigned( 162, 8)),
4 => std_logic_vector(to_unsigned( 148, 8)),
5 => std_logic_vector(to_unsigned( 113, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 111, 8)),
8 => std_logic_vector(to_unsigned( 93, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 88, 8)),
11 => std_logic_vector(to_unsigned( 109, 8)),
12 => std_logic_vector(to_unsigned( 91, 8)),
13 => std_logic_vector(to_unsigned( 119, 8)),
14 => std_logic_vector(to_unsigned( 115, 8)),
15 => std_logic_vector(to_unsigned( 67, 8)),
16 => std_logic_vector(to_unsigned( 91, 8)),
17 => std_logic_vector(to_unsigned( 88, 8)),
18 => std_logic_vector(to_unsigned( 108, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11101100
elsif count = 991 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 164, 8)),
2 => std_logic_vector(to_unsigned( 59, 8)),
3 => std_logic_vector(to_unsigned( 65, 8)),
4 => std_logic_vector(to_unsigned( 42, 8)),
5 => std_logic_vector(to_unsigned( 222, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 110, 8)),
8 => std_logic_vector(to_unsigned( 5, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 61, 8)),
11 => std_logic_vector(to_unsigned( 195, 8)),
12 => std_logic_vector(to_unsigned( 219, 8)),
13 => std_logic_vector(to_unsigned( 96, 8)),
14 => std_logic_vector(to_unsigned( 107, 8)),
15 => std_logic_vector(to_unsigned( 135, 8)),
16 => std_logic_vector(to_unsigned( 88, 8)),
17 => std_logic_vector(to_unsigned( 106, 8)),
18 => std_logic_vector(to_unsigned( 59, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011011
elsif count = 992 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 82, 8)),
2 => std_logic_vector(to_unsigned( 155, 8)),
3 => std_logic_vector(to_unsigned( 81, 8)),
4 => std_logic_vector(to_unsigned( 156, 8)),
5 => std_logic_vector(to_unsigned( 29, 8)),
6 => std_logic_vector(to_unsigned( 80, 8)),
7 => std_logic_vector(to_unsigned( 42, 8)),
8 => std_logic_vector(to_unsigned( 189, 8)),
9 => std_logic_vector(to_unsigned( 154, 8)),
10 => std_logic_vector(to_unsigned( 105, 8)),
11 => std_logic_vector(to_unsigned( 134, 8)),
12 => std_logic_vector(to_unsigned( 233, 8)),
13 => std_logic_vector(to_unsigned( 171, 8)),
14 => std_logic_vector(to_unsigned( 122, 8)),
15 => std_logic_vector(to_unsigned( 184, 8)),
16 => std_logic_vector(to_unsigned( 201, 8)),
17 => std_logic_vector(to_unsigned( 143, 8)),
18 => std_logic_vector(to_unsigned( 168, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11110011
elsif count = 993 then RAM <= (0 => "11111011",
1 => std_logic_vector(to_unsigned( 47, 8)),
2 => std_logic_vector(to_unsigned( 159, 8)),
3 => std_logic_vector(to_unsigned( 152, 8)),
4 => std_logic_vector(to_unsigned( 239, 8)),
5 => std_logic_vector(to_unsigned( 85, 8)),
6 => std_logic_vector(to_unsigned( 233, 8)),
7 => std_logic_vector(to_unsigned( 255, 8)),
8 => std_logic_vector(to_unsigned( 99, 8)),
9 => std_logic_vector(to_unsigned( 8, 8)),
10 => std_logic_vector(to_unsigned( 115, 8)),
11 => std_logic_vector(to_unsigned( 82, 8)),
12 => std_logic_vector(to_unsigned( 222, 8)),
13 => std_logic_vector(to_unsigned( 111, 8)),
14 => std_logic_vector(to_unsigned( 185, 8)),
15 => std_logic_vector(to_unsigned( 18, 8)),
16 => std_logic_vector(to_unsigned( 188, 8)),
17 => std_logic_vector(to_unsigned( 66, 8)),
18 => std_logic_vector(to_unsigned( 189, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11100001
elsif count = 994 then RAM <= (0 => "11111101",
1 => std_logic_vector(to_unsigned( 160, 8)),
2 => std_logic_vector(to_unsigned( 119, 8)),
3 => std_logic_vector(to_unsigned( 245, 8)),
4 => std_logic_vector(to_unsigned( 145, 8)),
5 => std_logic_vector(to_unsigned( 110, 8)),
6 => std_logic_vector(to_unsigned( 135, 8)),
7 => std_logic_vector(to_unsigned( 102, 8)),
8 => std_logic_vector(to_unsigned( 127, 8)),
9 => std_logic_vector(to_unsigned( 11, 8)),
10 => std_logic_vector(to_unsigned( 219, 8)),
11 => std_logic_vector(to_unsigned( 24, 8)),
12 => std_logic_vector(to_unsigned( 251, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 108, 8)),
15 => std_logic_vector(to_unsigned( 124, 8)),
16 => std_logic_vector(to_unsigned( 77, 8)),
17 => std_logic_vector(to_unsigned( 127, 8)),
18 => std_logic_vector(to_unsigned( 113, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11001101
elsif count = 995 then RAM <= (0 => "11110111",
1 => std_logic_vector(to_unsigned( 90, 8)),
2 => std_logic_vector(to_unsigned( 68, 8)),
3 => std_logic_vector(to_unsigned( 84, 8)),
4 => std_logic_vector(to_unsigned( 206, 8)),
5 => std_logic_vector(to_unsigned( 64, 8)),
6 => std_logic_vector(to_unsigned( 186, 8)),
7 => std_logic_vector(to_unsigned( 95, 8)),
8 => std_logic_vector(to_unsigned( 215, 8)),
9 => std_logic_vector(to_unsigned( 50, 8)),
10 => std_logic_vector(to_unsigned( 1, 8)),
11 => std_logic_vector(to_unsigned( 77, 8)),
12 => std_logic_vector(to_unsigned( 81, 8)),
13 => std_logic_vector(to_unsigned( 126, 8)),
14 => std_logic_vector(to_unsigned( 197, 8)),
15 => std_logic_vector(to_unsigned( 82, 8)),
16 => std_logic_vector(to_unsigned( 76, 8)),
17 => std_logic_vector(to_unsigned( 92, 8)),
18 => std_logic_vector(to_unsigned( 140, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10100111
elsif count = 996 then RAM <= (0 => "00111111",
1 => std_logic_vector(to_unsigned( 52, 8)),
2 => std_logic_vector(to_unsigned( 73, 8)),
3 => std_logic_vector(to_unsigned( 202, 8)),
4 => std_logic_vector(to_unsigned( 67, 8)),
5 => std_logic_vector(to_unsigned( 106, 8)),
6 => std_logic_vector(to_unsigned( 121, 8)),
7 => std_logic_vector(to_unsigned( 48, 8)),
8 => std_logic_vector(to_unsigned( 169, 8)),
9 => std_logic_vector(to_unsigned( 55, 8)),
10 => std_logic_vector(to_unsigned( 70, 8)),
11 => std_logic_vector(to_unsigned( 63, 8)),
12 => std_logic_vector(to_unsigned( 78, 8)),
13 => std_logic_vector(to_unsigned( 161, 8)),
14 => std_logic_vector(to_unsigned( 228, 8)),
15 => std_logic_vector(to_unsigned( 193, 8)),
16 => std_logic_vector(to_unsigned( 16, 8)),
17 => std_logic_vector(to_unsigned( 55, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 00111101
elsif count = 997 then RAM <= (0 => "10110111",
1 => std_logic_vector(to_unsigned( 83, 8)),
2 => std_logic_vector(to_unsigned( 59, 8)),
3 => std_logic_vector(to_unsigned( 102, 8)),
4 => std_logic_vector(to_unsigned( 110, 8)),
5 => std_logic_vector(to_unsigned( 127, 8)),
6 => std_logic_vector(to_unsigned( 133, 8)),
7 => std_logic_vector(to_unsigned( 199, 8)),
8 => std_logic_vector(to_unsigned( 226, 8)),
9 => std_logic_vector(to_unsigned( 208, 8)),
10 => std_logic_vector(to_unsigned( 70, 8)),
11 => std_logic_vector(to_unsigned( 178, 8)),
12 => std_logic_vector(to_unsigned( 40, 8)),
13 => std_logic_vector(to_unsigned( 151, 8)),
14 => std_logic_vector(to_unsigned( 18, 8)),
15 => std_logic_vector(to_unsigned( 206, 8)),
16 => std_logic_vector(to_unsigned( 124, 8)),
17 => std_logic_vector(to_unsigned( 162, 8)),
18 => std_logic_vector(to_unsigned( 96, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 10110100
elsif count = 998 then RAM <= (0 => "11011011",
1 => std_logic_vector(to_unsigned( 249, 8)),
2 => std_logic_vector(to_unsigned( 113, 8)),
3 => std_logic_vector(to_unsigned( 147, 8)),
4 => std_logic_vector(to_unsigned( 155, 8)),
5 => std_logic_vector(to_unsigned( 199, 8)),
6 => std_logic_vector(to_unsigned( 226, 8)),
7 => std_logic_vector(to_unsigned( 174, 8)),
8 => std_logic_vector(to_unsigned( 64, 8)),
9 => std_logic_vector(to_unsigned( 219, 8)),
10 => std_logic_vector(to_unsigned( 143, 8)),
11 => std_logic_vector(to_unsigned( 184, 8)),
12 => std_logic_vector(to_unsigned( 68, 8)),
13 => std_logic_vector(to_unsigned( 147, 8)),
14 => std_logic_vector(to_unsigned( 155, 8)),
15 => std_logic_vector(to_unsigned( 145, 8)),
16 => std_logic_vector(to_unsigned( 153, 8)),
17 => std_logic_vector(to_unsigned( 177, 8)),
18 => std_logic_vector(to_unsigned( 123, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 11011010
elsif count = 999 then RAM <= (0 => "11110110",
1 => std_logic_vector(to_unsigned( 138, 8)),
2 => std_logic_vector(to_unsigned( 2, 8)),
3 => std_logic_vector(to_unsigned( 176, 8)),
4 => std_logic_vector(to_unsigned( 53, 8)),
5 => std_logic_vector(to_unsigned( 71, 8)),
6 => std_logic_vector(to_unsigned( 191, 8)),
7 => std_logic_vector(to_unsigned( 158, 8)),
8 => std_logic_vector(to_unsigned( 150, 8)),
9 => std_logic_vector(to_unsigned( 140, 8)),
10 => std_logic_vector(to_unsigned( 113, 8)),
11 => std_logic_vector(to_unsigned( 171, 8)),
12 => std_logic_vector(to_unsigned( 144, 8)),
13 => std_logic_vector(to_unsigned( 133, 8)),
14 => std_logic_vector(to_unsigned( 106, 8)),
15 => std_logic_vector(to_unsigned( 119, 8)),
16 => std_logic_vector(to_unsigned( 8, 8)),
17 => std_logic_vector(to_unsigned( 190, 8)),
18 => std_logic_vector(to_unsigned( 101, 8)),
 others => (others => '0'));
-- MASK_OUT: 	 01110010
end if; end if;
                end process;
                test : process is
                begin  wait for 100 ns;
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '1';
                    wait for c_CLOCK_PERIOD;
                    tb_rst <= '0';   wait for c_CLOCK_PERIOD;
                    count <= 0;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 1;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 2;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 3;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 4;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 5;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 6;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 7;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 8;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 9;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 10;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 11;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 12;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 13;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 14;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 15;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 16;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 17;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 18;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 19;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 20;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 21;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 22;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 23;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 24;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 25;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 26;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 27;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 28;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 29;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 30;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 31;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 32;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 33;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 34;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 35;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 36;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 37;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 38;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 39;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 40;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 41;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 42;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 43;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 44;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 45;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 46;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 47;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 48;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 49;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 50;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 51;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 52;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 53;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 54;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 55;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 56;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 57;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 58;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 59;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 60;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 61;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 62;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 63;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 64;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 65;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 66;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 67;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 68;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 69;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 70;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 71;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 72;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 73;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 74;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 75;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 76;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 77;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 78;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 79;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 80;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 81;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 82;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 83;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 84;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 85;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 86;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 87;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 88;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 89;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 90;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 91;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 92;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 93;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 94;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 95;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 96;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 97;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 98;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 99;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 100;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 101;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 102;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 103;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 104;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 105;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 106;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 107;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 108;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 109;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 110;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 111;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 112;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 113;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 114;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 115;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 116;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 117;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 118;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 119;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 120;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 121;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 122;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 123;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 124;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 125;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 126;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 127;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 128;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 129;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 130;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 131;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 132;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 133;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 134;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 135;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 136;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 137;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 138;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 139;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 140;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 141;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 142;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 143;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 144;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 145;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 146;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 147;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 148;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 149;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 150;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 151;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 152;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 153;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 154;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 155;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 156;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 157;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 158;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 159;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 160;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 161;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 162;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 163;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 164;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 165;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 166;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 167;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 168;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 169;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 170;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 171;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 172;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 173;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 174;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 175;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 176;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 177;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 178;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 179;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 180;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 181;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 182;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 183;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 184;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 185;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 186;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 187;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 188;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 189;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 190;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 191;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 192;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 193;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 194;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 195;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 196;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 197;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 198;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 199;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 200;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 201;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 202;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 203;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 204;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 205;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 206;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 207;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 208;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 209;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 210;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 211;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 212;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 213;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 214;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 215;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 216;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 217;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 218;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 219;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 220;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 221;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 222;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 223;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 224;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 225;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 226;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 227;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 228;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 229;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 230;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 231;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 232;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 233;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 234;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 235;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 236;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 237;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 238;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 239;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 240;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 241;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 242;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 243;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 244;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 245;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 246;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 247;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 248;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 249;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 250;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 251;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 252;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 253;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 254;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 255;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 256;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 257;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 258;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 259;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 260;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 261;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 262;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 263;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 264;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 265;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 266;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 267;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 268;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 269;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 270;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 271;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 272;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 273;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 274;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 275;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 276;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 277;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 278;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 279;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 280;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 281;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 282;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 283;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 284;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 285;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 286;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 287;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 288;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 289;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 290;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 291;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 292;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 293;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 294;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 295;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 296;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 297;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 298;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 299;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 300;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 301;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 302;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 303;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 304;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 305;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 306;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 307;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 308;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 309;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 310;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 311;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 312;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 313;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 314;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 315;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 316;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 317;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 318;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 319;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 320;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 321;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 322;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 323;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 324;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 325;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 326;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 327;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 328;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 329;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 330;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 331;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 332;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 333;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 334;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 335;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 336;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 337;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 338;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 339;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 340;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 341;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 342;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 343;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 344;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 345;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 346;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 347;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 348;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 349;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 350;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 351;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 352;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 353;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 354;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 355;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 356;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 357;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 358;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 359;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 360;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 361;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 362;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 363;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 364;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 365;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 366;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 367;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 368;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 369;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 370;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 371;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 372;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 373;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 374;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 375;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 376;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 377;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 378;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 379;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 380;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 381;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 382;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 383;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 384;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 385;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 386;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 387;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 388;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 389;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 390;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 391;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 392;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 393;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 394;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 395;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 396;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 397;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 398;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 399;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 400;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 401;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 402;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 403;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 404;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 405;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 406;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 407;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 408;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 409;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 410;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 411;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 412;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 413;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 414;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 415;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 416;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 417;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 418;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 419;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 420;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 421;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 422;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 423;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 424;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 425;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 426;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 427;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 428;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 429;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 430;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 431;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 432;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 433;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 434;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 435;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 436;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 437;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 438;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 439;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 440;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 441;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 442;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 443;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 444;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 445;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 446;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 447;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 448;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 449;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 450;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 451;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 452;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 453;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 454;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 455;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 456;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 457;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 458;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 459;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 460;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 461;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 462;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 463;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 464;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 465;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 466;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 467;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 468;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 469;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 470;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 471;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 472;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 473;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 474;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 475;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 476;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 477;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 478;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 479;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 480;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 481;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 482;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 483;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 484;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 485;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 486;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 487;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 488;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 489;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 490;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 491;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 492;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 493;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 494;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 495;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 496;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 497;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 498;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 499;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 500;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 501;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 502;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 503;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 504;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 505;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 506;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 507;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 508;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 509;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 510;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 511;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 512;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 513;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 514;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 515;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 516;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 517;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 518;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 519;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 520;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 521;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 522;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 523;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 524;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 525;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 526;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 527;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 528;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 529;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 530;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 531;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 532;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 533;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 534;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 535;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 536;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 537;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 538;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 539;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 540;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 541;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 542;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 543;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 544;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 545;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 546;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 547;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 548;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 549;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 550;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 551;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 552;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 553;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 554;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 555;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 556;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 557;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 558;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 559;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 560;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 561;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 562;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 563;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 564;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 565;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 566;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 567;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 568;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 569;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 570;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 571;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 572;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 573;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 574;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 575;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 576;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 577;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 578;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 579;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 580;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 581;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 582;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 583;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 584;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 585;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 586;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 587;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 588;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 589;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 590;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 591;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 592;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 593;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 594;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 595;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 596;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 597;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 598;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 599;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 600;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 601;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 602;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 603;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 604;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 605;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 606;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 607;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 608;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 609;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 610;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 611;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 612;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 613;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 614;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 615;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 616;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 617;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 618;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 619;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 620;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 621;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 622;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 623;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 624;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 625;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 626;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 627;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 628;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 629;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 630;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 631;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 632;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 633;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 634;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 635;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 636;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 637;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 638;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 639;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 640;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 641;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 642;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 643;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 644;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 645;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 646;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 647;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 648;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 649;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 650;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 651;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 652;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 653;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 654;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 655;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 656;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 657;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 658;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 659;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 660;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 661;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 662;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 663;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 664;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 665;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 666;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 667;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 668;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 669;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 670;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 671;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 672;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 673;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 674;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 675;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 676;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 677;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 678;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 679;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 680;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 681;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 682;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 683;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 684;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 685;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 686;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 687;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 688;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 689;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 690;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 691;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 692;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 693;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 694;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 695;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 696;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 697;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 698;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 699;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 700;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 701;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 702;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 703;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 704;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 705;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 706;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 707;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 708;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 709;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 710;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 711;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 712;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 713;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 714;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 715;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 716;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 717;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 718;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 719;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 720;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 721;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 722;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 723;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 724;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 725;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 726;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 727;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 728;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 729;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 730;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 731;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 732;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 733;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 734;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 735;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 736;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 737;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 738;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 739;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 740;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 741;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 742;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 743;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 744;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 745;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 746;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 747;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 748;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 749;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 750;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 751;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 752;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 753;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 754;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 755;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 756;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 757;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 758;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 759;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 760;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 761;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 762;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 763;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 764;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 765;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 766;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 767;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 768;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 769;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 770;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 771;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 772;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 773;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 774;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 775;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 776;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 777;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 778;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 779;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 780;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 781;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 782;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 783;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 784;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 785;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 786;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 787;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 788;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 789;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 790;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 791;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 792;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 793;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 794;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 795;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 796;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 797;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 798;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 799;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 800;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 801;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 802;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 803;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 804;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 805;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 806;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 807;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 808;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 809;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 810;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 811;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 812;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 813;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 814;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 815;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 816;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 817;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 818;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 819;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 820;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 821;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 822;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 823;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 824;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 825;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 826;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 827;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 828;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 829;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 830;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 831;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 832;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 833;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 834;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 835;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 836;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 837;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 838;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 839;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 840;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 841;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 842;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 843;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 844;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 845;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 846;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 847;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 848;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 849;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 850;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 851;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 852;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 853;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 854;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 855;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 856;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 857;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 858;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 859;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 860;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 861;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 862;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 863;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 864;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 865;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 866;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 867;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 868;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 869;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 870;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 871;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 872;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 873;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 874;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 875;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 876;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 877;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 878;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 879;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 880;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 881;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 882;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 883;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 884;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 885;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 886;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 887;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 888;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 889;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 890;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 891;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 892;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 893;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 894;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 895;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 896;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 897;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 898;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 899;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 900;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 901;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 902;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 903;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 904;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 905;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 906;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 907;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 908;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 909;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 910;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 911;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10000111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 912;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 913;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 914;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 915;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 916;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 917;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 918;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 919;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 920;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 921;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110000" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 922;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 923;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 924;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 925;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 926;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 927;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 928;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 929;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 930;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 931;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 932;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 933;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 934;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 935;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 936;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 937;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 938;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 939;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 940;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 941;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 942;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11010010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 943;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00110110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 944;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 945;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 946;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 947;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 948;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 949;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 950;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 951;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 952;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 953;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 954;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 955;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 956;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11000011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 957;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 958;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 959;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10111110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 960;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 961;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01001011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 962;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 963;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 964;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 965;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 966;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 967;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 968;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 969;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 970;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01111011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 971;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 972;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 973;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 974;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 975;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00101111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 976;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 977;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10011111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 978;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 979;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 980;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 981;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00010111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 982;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00011110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 983;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 984;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10101010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 985;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 986;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 987;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 988;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11111010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 989;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01010110" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 990;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11101100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 991;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 992;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11110011" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 993;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11100001" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 994;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11001101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 995;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10100111" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 996;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "00111101" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 997;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "10110100" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 998;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "11011010" report "TEST FAILED" severity failure;  wait for c_CLOCK_PERIOD;
                    count <= 999;
                    wait for c_CLOCK_PERIOD;
                    count <= 0;
                    tb_start <= '1';
                    wait for c_CLOCK_PERIOD;
                    wait until tb_done = '1';
                    wait for c_CLOCK_PERIOD;
                    tb_start <= '0';
                    wait until tb_done = '0';
                    assert RAM(19) = "01110010" report "TEST FAILED" severity failure;
assert false report "1000 TESTS PASSED" severity failure;
    end process test;
                end projecttb;